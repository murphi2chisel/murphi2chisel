module Store(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h1 : io_Sta_in_Proc_1_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h1 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h2 : io_Sta_in_Proc_1_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h2 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h1 : io_Sta_in_Proc_2_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h1 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h2 : io_Sta_in_Proc_2_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h2 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_4(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h1 : io_Sta_in_Proc_3_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h1 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h2 : io_Sta_in_Proc_3_CacheData; // @[router.scala 13:49 14:32 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h2 : io_Sta_in_CurrData; // @[router.scala 13:49 15:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheData; // @[router.scala 12:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 12:14 node.scala 25:11]
endmodule
module Store_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeProc_CacheState == 2'h2 ? 2'h1 : io_Sta_in_HomeProc_CacheData; // @[router.scala 21:48 22:31 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_HomeProc_CacheState == 2'h2 ? 2'h1 : io_Sta_in_CurrData; // @[router.scala 21:48 23:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_en_r ? _GEN_0 : io_Sta_in_HomeProc_CacheData; // @[router.scala 20:14 node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 20:14 node.scala 25:11]
endmodule
module Store_Home_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeProc_CacheState == 2'h2 ? 2'h2 : io_Sta_in_HomeProc_CacheData; // @[router.scala 21:48 22:31 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_HomeProc_CacheState == 2'h2 ? 2'h2 : io_Sta_in_CurrData; // @[router.scala 21:48 23:21 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_en_r ? _GEN_0 : io_Sta_in_HomeProc_CacheData; // @[router.scala 20:14 node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_en_r ? _GEN_1 : io_Sta_in_CurrData; // @[router.scala 20:14 node.scala 25:11]
endmodule
module PI_Remote_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 ? 2'h1 :
    io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11 router.scala 29:94 30:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 ? 3'h1 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 29:94 31:28]
  wire  _GEN_2 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 | io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 29:94 32:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_Get_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 ? 2'h1 :
    io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11 router.scala 29:94 30:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 ? 3'h1 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 29:94 31:28]
  wire  _GEN_2 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 | io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 29:94 32:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_Get_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 ? 2'h1 :
    io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11 router.scala 29:94 30:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 ? 3'h1 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 29:94 31:28]
  wire  _GEN_2 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 | io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 29:94 32:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 28:14]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_Get_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~
    io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? 2'h1 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 38:143 39:29]
  wire  _GEN_1 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~io_Sta_in_Dir_Pending
     & io_Sta_in_Dir_Dirty)) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 38:143 40:24]
  wire [2:0] _GEN_2 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~
    io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? 3'h1 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 38:143 41:27]
  wire [1:0] _GEN_3 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~
    io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? io_Sta_in_Dir_HeadPtr : io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11 router.scala 38:143 42:28]
  wire  _GEN_4 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~io_Sta_in_Dir_Pending
     & io_Sta_in_Dir_Dirty)) ? io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11 router.scala 38:143 43:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 37:14]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_1 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 37:14]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_2 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 37:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_en_r ? _GEN_3 : io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11 router.scala 37:14]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_en_r ? _GEN_4 : io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11 router.scala 37:14]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_Get_Put(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_HomeProc_InvMarked ? 1'h0 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 52:35 53:31]
  wire  _GEN_1 = io_Sta_in_HomeProc_InvMarked ? 1'h0 : 1'h1; // @[router.scala 52:35 54:32 56:32]
  wire  _GEN_2 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~io_Sta_in_Dir_Pending
     & ~io_Sta_in_Dir_Dirty)) | io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 49:146 50:22]
  wire [1:0] _GEN_3 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~
    io_Sta_in_Dir_Pending & ~io_Sta_in_Dir_Dirty)) ? 2'h0 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 49:146 51:29]
  wire  _GEN_4 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~io_Sta_in_Dir_Pending
     & ~io_Sta_in_Dir_Dirty)) ? _GEN_0 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 49:146]
  wire [1:0] _GEN_5 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & (io_Sta_in_HomeProc_CacheState == 2'h0 & (~
    io_Sta_in_Dir_Pending & ~io_Sta_in_Dir_Dirty)) ? {{1'd0}, _GEN_1} : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 49:146]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_3 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 48:14]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_4 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 48:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_5 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 48:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_2 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 48:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_GetX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 ? 2'h2 :
    io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11 router.scala 64:94 65:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 ? 3'h2 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 64:94 66:28]
  wire  _GEN_2 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h0 | io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 64:94 67:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_GetX_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 ? 2'h2 :
    io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11 router.scala 64:94 65:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 ? 3'h2 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 64:94 66:28]
  wire  _GEN_2 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h0 | io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 64:94 67:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_GetX_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 ? 2'h2 :
    io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11 router.scala 64:94 65:30]
  wire [2:0] _GEN_1 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 ? 3'h2 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 64:94 66:28]
  wire  _GEN_2 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h0 | io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 64:94 67:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 63:14]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_GetX_GetX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? 2'h2 :
    io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 73:188 74:29]
  wire  _GEN_1 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 73:188 75:24]
  wire [2:0] _GEN_2 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? 3'h2 :
    io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 73:188 76:27]
  wire [1:0] _GEN_3 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? io_Sta_in_Dir_HeadPtr :
    io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11 router.scala 73:188 77:28]
  wire  _GEN_4 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & io_Sta_in_Dir_Dirty)) ? io_Sta_in_Dir_HomeHeadPtr
     : io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11 router.scala 73:188 78:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_0 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 72:14]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_1 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 72:14]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_2 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 72:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_en_r ? _GEN_3 : io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11 router.scala 72:14]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_en_r ? _GEN_4 : io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11 router.scala 72:14]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_GetX_PutX_HeadVld(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_14 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadPtr == 2'h1 & ~
    io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 92:54]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadPtr == 2'h1 & ~
    io_Sta_in_Dir_HomeHeadPtr ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 92:119 94:26]
  wire  _T_19 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadPtr == 2'h2 & ~
    io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 92:54]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadPtr == 2'h2 & ~
    io_Sta_in_Dir_HomeHeadPtr ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 92:119 94:26]
  wire  _T_24 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadPtr == 2'h3 & ~
    io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 92:54]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadPtr == 2'h3 & ~
    io_Sta_in_Dir_HomeHeadPtr ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 92:119 94:26]
  wire  _GEN_6 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     | io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 84:216 85:22]
  wire  _GEN_7 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 84:216 86:22]
  wire  _GEN_8 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 84:216 87:24]
  wire  _GEN_9 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 84:216 88:24]
  wire  _GEN_10 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 84:216 89:23]
  wire  _GEN_11 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 84:216 91:26]
  wire  _GEN_12 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _T_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 84:216]
  wire [1:0] _GEN_13 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 84:216]
  wire  _GEN_14 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 84:216 91:26]
  wire  _GEN_15 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _T_19 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 84:216]
  wire [1:0] _GEN_16 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 84:216]
  wire  _GEN_17 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 84:216 91:26]
  wire  _GEN_18 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _T_24 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 84:216]
  wire [1:0] _GEN_19 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 84:216]
  wire  _GEN_20 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[router.scala 84:216 101:27 node.scala 25:11]
  wire  _GEN_21 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[router.scala 84:216 102:27 node.scala 25:11]
  wire [1:0] _GEN_22 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[router.scala 84:216 103:27 node.scala 25:11]
  wire [1:0] _GEN_23 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 2'h0 : io_Sta_in_HomeProc_ProcCmd; // @[router.scala 84:216 104:29 node.scala 25:11]
  wire  _GEN_24 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_HomeProc_InvMarked; // @[router.scala 84:216 105:31 node.scala 25:11]
  wire [1:0] _GEN_25 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? 2'h2 : io_Sta_in_HomeProc_CacheState; // @[router.scala 84:216 106:32 node.scala 25:11]
  wire [1:0] _GEN_26 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))
     ? io_Sta_in_MemData : io_Sta_in_HomeProc_CacheData; // @[router.scala 84:216 107:31 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_23 : io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_24 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_25 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_HomeProc_CacheData = io_en_r ? _GEN_26 : io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_8 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_6 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_7 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_11 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_14 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_17 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_20 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_12 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_15 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_18 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_21 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_13 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_16 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_19 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_22 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 83:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_GetX_PutX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     | io_Sta_in_Dir_Local; // @[router.scala 113:219 114:22 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     | io_Sta_in_Dir_Dirty; // @[router.scala 113:219 115:22 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     ? 2'h0 : io_Sta_in_HomeProc_ProcCmd; // @[router.scala 113:219 116:29 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     ? 1'h0 : io_Sta_in_HomeProc_InvMarked; // @[router.scala 113:219 117:31 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     ? 2'h2 : io_Sta_in_HomeProc_CacheState; // @[router.scala 113:219 118:32 node.scala 25:11]
  wire [1:0] _GEN_5 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & ((io_Sta_in_HomeProc_CacheState == 2'h0 |
    io_Sta_in_HomeProc_CacheState == 2'h1) & (~io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))
     ? io_Sta_in_MemData : io_Sta_in_HomeProc_CacheData; // @[router.scala 113:219 119:31 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_2 : io_Sta_in_HomeProc_ProcCmd; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_3 : io_Sta_in_HomeProc_InvMarked; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_4 : io_Sta_in_HomeProc_CacheState; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_en_r ? _GEN_5 : io_Sta_in_HomeProc_CacheData; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[router.scala 112:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_PutX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h0 :
    io_Sta_in_Proc_1_CacheState; // @[router.scala 125:94 126:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h2 | io_Sta_in_WbMsg_Cmd; // @[router.scala 125:94 127:22 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h2 ? 2'h1 :
    io_Sta_in_WbMsg_Proc; // @[router.scala 125:94 128:23 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h2 ? 1'h0 :
    io_Sta_in_WbMsg_HomeProc; // @[router.scala 125:94 129:27 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h2 ?
    io_Sta_in_Proc_1_CacheData : io_Sta_in_WbMsg_Data; // @[router.scala 125:94 130:23 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheState; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_WbMsg_Cmd; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_en_r ? _GEN_2 : io_Sta_in_WbMsg_Proc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_WbMsg_HomeProc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_en_r ? _GEN_4 : io_Sta_in_WbMsg_Data; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_PutX_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h0 :
    io_Sta_in_Proc_2_CacheState; // @[router.scala 125:94 126:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h2 | io_Sta_in_WbMsg_Cmd; // @[router.scala 125:94 127:22 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h2 ? 2'h2 :
    io_Sta_in_WbMsg_Proc; // @[router.scala 125:94 128:23 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h2 ? 1'h0 :
    io_Sta_in_WbMsg_HomeProc; // @[router.scala 125:94 129:27 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h2 ?
    io_Sta_in_Proc_2_CacheData : io_Sta_in_WbMsg_Data; // @[router.scala 125:94 130:23 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheState; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_WbMsg_Cmd; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_en_r ? _GEN_2 : io_Sta_in_WbMsg_Proc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_WbMsg_HomeProc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_en_r ? _GEN_4 : io_Sta_in_WbMsg_Data; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_PutX_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h0 :
    io_Sta_in_Proc_3_CacheState; // @[router.scala 125:94 126:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h2 | io_Sta_in_WbMsg_Cmd; // @[router.scala 125:94 127:22 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h2 ? 2'h3 :
    io_Sta_in_WbMsg_Proc; // @[router.scala 125:94 128:23 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h2 ? 1'h0 :
    io_Sta_in_WbMsg_HomeProc; // @[router.scala 125:94 129:27 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h2 ?
    io_Sta_in_Proc_3_CacheData : io_Sta_in_WbMsg_Data; // @[router.scala 125:94 130:23 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheState; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_WbMsg_Cmd; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_en_r ? _GEN_2 : io_Sta_in_WbMsg_Proc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_WbMsg_HomeProc; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_en_r ? _GEN_4 : io_Sta_in_WbMsg_Data; // @[router.scala 124:14 node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_PutX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_1 = io_Sta_in_Dir_Pending ? 1'h0 : io_Sta_in_Dir_Dirty; // @[router.scala 137:28 139:22 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_Dir_Pending ? io_Sta_in_HomeProc_CacheData : io_Sta_in_MemData; // @[router.scala 137:28 140:20 node.scala 25:11]
  wire [1:0] _GEN_3 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & io_Sta_in_HomeProc_CacheState == 2'h2 ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[router.scala 136:92 node.scala 25:11]
  wire  _GEN_4 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & io_Sta_in_HomeProc_CacheState == 2'h2 ? _GEN_1 :
    io_Sta_in_Dir_Dirty; // @[router.scala 136:92 node.scala 25:11]
  wire [1:0] _GEN_5 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & io_Sta_in_HomeProc_CacheState == 2'h2 ? _GEN_2 :
    io_Sta_in_MemData; // @[router.scala 136:92 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_3 : io_Sta_in_HomeProc_CacheState; // @[router.scala 135:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_4 : io_Sta_in_Dir_Dirty; // @[router.scala 135:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_en_r ? _GEN_5 : io_Sta_in_MemData; // @[router.scala 135:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_Replace(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h1 ? 2'h0 :
    io_Sta_in_Proc_1_CacheState; // @[router.scala 150:94 151:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_1_ProcCmd == 2'h0 & io_Sta_in_Proc_1_CacheState == 2'h1 | io_Sta_in_RpMsg_1_Cmd; // @[router.scala 150:94 152:27 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheState; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_RpMsg_1_Cmd; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_Replace_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h1 ? 2'h0 :
    io_Sta_in_Proc_2_CacheState; // @[router.scala 150:94 151:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_2_ProcCmd == 2'h0 & io_Sta_in_Proc_2_CacheState == 2'h1 | io_Sta_in_RpMsg_2_Cmd; // @[router.scala 150:94 152:27 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheState; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_RpMsg_2_Cmd; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Remote_Replace_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h1 ? 2'h0 :
    io_Sta_in_Proc_3_CacheState; // @[router.scala 150:94 151:33 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_Proc_3_ProcCmd == 2'h0 & io_Sta_in_Proc_3_CacheState == 2'h1 | io_Sta_in_RpMsg_3_Cmd; // @[router.scala 150:94 152:27 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheState; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_RpMsg_3_Cmd; // @[router.scala 149:14 node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module PI_Local_Replace(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & io_Sta_in_HomeProc_CacheState == 2'h1 ? 1'h0 : io_Sta_in_Dir_Local
    ; // @[router.scala 158:92 159:22 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_HomeProc_ProcCmd == 2'h0 & io_Sta_in_HomeProc_CacheState == 2'h1 ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[router.scala 158:92 160:32 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_1 : io_Sta_in_HomeProc_CacheState; // @[router.scala 157:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[router.scala 157:14 node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Nak(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h5 ? 3'h0 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 166:44 167:28 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h5 ? 2'h0 : io_Sta_in_Proc_1_ProcCmd; // @[router.scala 166:44 168:30 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h5 ? 1'h0 : io_Sta_in_Proc_1_InvMarked; // @[router.scala 166:44 169:32 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_en_r ? _GEN_1 : io_Sta_in_Proc_1_ProcCmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_en_r ? _GEN_2 : io_Sta_in_Proc_1_InvMarked; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Nak_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h5 ? 3'h0 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 166:44 167:28 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h5 ? 2'h0 : io_Sta_in_Proc_2_ProcCmd; // @[router.scala 166:44 168:30 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h5 ? 1'h0 : io_Sta_in_Proc_2_InvMarked; // @[router.scala 166:44 169:32 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_en_r ? _GEN_1 : io_Sta_in_Proc_2_ProcCmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_en_r ? _GEN_2 : io_Sta_in_Proc_2_InvMarked; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Nak_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h5 ? 3'h0 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 166:44 167:28 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h5 ? 2'h0 : io_Sta_in_Proc_3_ProcCmd; // @[router.scala 166:44 168:30 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h5 ? 1'h0 : io_Sta_in_Proc_3_InvMarked; // @[router.scala 166:44 169:32 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_en_r ? _GEN_1 : io_Sta_in_Proc_3_ProcCmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_en_r ? _GEN_2 : io_Sta_in_Proc_3_InvMarked; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 165:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Nak_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h5 ? 3'h0 : io_Sta_in_HomeUniMsg_Cmd; // @[router.scala 175:43 176:27 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h5 ? 2'h0 : io_Sta_in_HomeProc_ProcCmd; // @[router.scala 175:43 177:29 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_HomeUniMsg_Cmd == 3'h5 ? 1'h0 : io_Sta_in_HomeProc_InvMarked; // @[router.scala 175:43 178:31 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_en_r ? _GEN_1 : io_Sta_in_HomeProc_ProcCmd; // @[router.scala 174:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_2 : io_Sta_in_HomeProc_InvMarked; // @[router.scala 174:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_0 : io_Sta_in_HomeUniMsg_Cmd; // @[router.scala 174:14 node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Nak_Clear(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_NakcMsg_Cmd ? 1'h0 : io_Sta_in_NakcMsg_Cmd; // @[router.scala 184:42 185:24 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_NakcMsg_Cmd ? 1'h0 : io_Sta_in_Dir_Pending; // @[router.scala 184:42 186:24 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_1 : io_Sta_in_Dir_Pending; // @[router.scala 183:14 node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_0 : io_Sta_in_NakcMsg_Cmd; // @[router.scala 183:14 node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Nak(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (
    io_Sta_in_Dir_Pending | (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) |
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h1 & ~io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h5
     : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 192:353 193:28 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 191:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Nak_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (
    io_Sta_in_Dir_Pending | (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) |
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h2 & ~io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h5
     : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 192:353 193:28 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 191:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Nak_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (
    io_Sta_in_Dir_Pending | (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) |
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h3 & ~io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h5
     : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 192:353 193:28 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 191:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 |
    io_Sta_in_Dir_HomeHeadPtr)))))) | io_Sta_in_Dir_Pending; // @[router.scala 199:262 200:24 node.scala 25:11]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h1 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 199:262 201:28 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_1_Proc; // @[router.scala 199:262 202:29 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_1_HomeProc; // @[router.scala 199:262 203:33 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_Proc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_1_HomeProc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Get_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 |
    io_Sta_in_Dir_HomeHeadPtr)))))) | io_Sta_in_Dir_Pending; // @[router.scala 199:262 200:24 node.scala 25:11]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h1 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 199:262 201:28 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_2_Proc; // @[router.scala 199:262 202:29 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_2_HomeProc; // @[router.scala 199:262 203:33 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_Proc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_2_HomeProc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Get_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 |
    io_Sta_in_Dir_HomeHeadPtr)))))) | io_Sta_in_Dir_Pending; // @[router.scala 199:262 200:24 node.scala 25:11]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? 3'h1 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 199:262 201:28 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_3_Proc; // @[router.scala 199:262 202:29 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 |
    io_Sta_in_Dir_HomeHeadPtr)))))) ? io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_3_HomeProc; // @[router.scala 199:262 203:33 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_Proc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_3_HomeProc; // @[router.scala 198:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Head(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrVld; // @[router.scala 209:200 210:23 node.scala 25:11]
  wire  _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrSet_1; // @[router.scala 209:200 211:28 node.scala 25:11]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_InvSet_1; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_2 :
    io_Sta_in_Dir_InvSet_2; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_3 :
    io_Sta_in_Dir_InvSet_3; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_HomeShrSet :
    io_Sta_in_Dir_HomeInvSet; // @[router.scala 209:200 221:27 node.scala 25:11]
  wire [2:0] _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 209:200 222:28 node.scala 25:11]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[router.scala 209:200 223:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_3 : io_Sta_in_Dir_ShrVld; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_4 : io_Sta_in_Dir_ShrSet_1; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_5 : io_Sta_in_Dir_InvSet_1; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_6 : io_Sta_in_Dir_InvSet_2; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_3; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_8 : io_Sta_in_Dir_HomeInvSet; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_9 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_10 : io_Sta_in_UniMsg_1_Data; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Head_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrVld; // @[router.scala 209:200 210:23 node.scala 25:11]
  wire  _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrSet_2; // @[router.scala 209:200 211:28 node.scala 25:11]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_1 :
    io_Sta_in_Dir_InvSet_1; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_InvSet_2; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_3 :
    io_Sta_in_Dir_InvSet_3; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_HomeShrSet :
    io_Sta_in_Dir_HomeInvSet; // @[router.scala 209:200 221:27 node.scala 25:11]
  wire [2:0] _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 209:200 222:28 node.scala 25:11]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[router.scala 209:200 223:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_3 : io_Sta_in_Dir_ShrVld; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_4 : io_Sta_in_Dir_ShrSet_2; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_5 : io_Sta_in_Dir_InvSet_1; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_6 : io_Sta_in_Dir_InvSet_2; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_3; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_8 : io_Sta_in_Dir_HomeInvSet; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_9 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_10 : io_Sta_in_UniMsg_2_Data; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Head_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrVld; // @[router.scala 209:200 210:23 node.scala 25:11]
  wire  _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_ShrSet_3; // @[router.scala 209:200 211:28 node.scala 25:11]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_1 :
    io_Sta_in_Dir_InvSet_1; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_ShrSet_2 :
    io_Sta_in_Dir_InvSet_2; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_InvSet_3; // @[router.scala 209:200 node.scala 25:11]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_Dir_HomeShrSet :
    io_Sta_in_Dir_HomeInvSet; // @[router.scala 209:200 221:27 node.scala 25:11]
  wire [2:0] _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 209:200 222:28 node.scala 25:11]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[router.scala 209:200 223:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_3 : io_Sta_in_Dir_ShrVld; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_4 : io_Sta_in_Dir_ShrSet_3; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_5 : io_Sta_in_Dir_InvSet_1; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_6 : io_Sta_in_Dir_InvSet_2; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_3; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_8 : io_Sta_in_Dir_HomeInvSet; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_9 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_10 : io_Sta_in_UniMsg_3_Data; // @[router.scala 208:14 node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_HeadVld; // @[router.scala 229:203 230:24 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[router.scala 229:203 231:24 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 229:203 232:28 node.scala 25:11]
  wire [2:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 229:203 233:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[router.scala 229:203 234:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_0 : io_Sta_in_Dir_HeadVld; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_4 : io_Sta_in_UniMsg_1_Data; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_HeadVld; // @[router.scala 229:203 230:24 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[router.scala 229:203 231:24 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 229:203 232:28 node.scala 25:11]
  wire [2:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 229:203 233:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[router.scala 229:203 234:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_0 : io_Sta_in_Dir_HeadVld; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_4 : io_Sta_in_UniMsg_2_Data; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) | io_Sta_in_Dir_HeadVld; // @[router.scala 229:203 230:24 node.scala 25:11]
  wire [1:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[router.scala 229:203 231:24 node.scala 25:11]
  wire  _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 229:203 232:28 node.scala 25:11]
  wire [2:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? 3'h3 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 229:203 233:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (~io_Sta_in_Dir_Dirty & ~io_Sta_in_Dir_HeadVld)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[router.scala 229:203 234:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_0 : io_Sta_in_Dir_HeadVld; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_4 : io_Sta_in_UniMsg_3_Data; // @[router.scala 228:14 node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Dirty(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_Dirty; // @[router.scala 240:240 241:22 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) |
    io_Sta_in_Dir_HeadVld; // @[router.scala 240:240 242:24 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h1
     : io_Sta_in_Dir_HeadPtr; // @[router.scala 240:240 243:24 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 240:240 244:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_MemData; // @[router.scala 240:240 245:20 node.scala 25:11]
  wire [1:0] _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h1
     : io_Sta_in_HomeProc_CacheState; // @[router.scala 240:240 246:32 node.scala 25:11]
  wire [2:0] _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 3'h3
     : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 240:240 247:28 node.scala 25:11]
  wire [1:0] _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_RpMsg_1_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_UniMsg_1_Data; // @[router.scala 240:240 248:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_5 : io_Sta_in_HomeProc_CacheState; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_0 : io_Sta_in_Dir_Dirty; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadVld; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_en_r ? _GEN_4 : io_Sta_in_MemData; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_6 : io_Sta_in_UniMsg_1_Cmd; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_7 : io_Sta_in_UniMsg_1_Data; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Dirty_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_Dirty; // @[router.scala 240:240 241:22 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) |
    io_Sta_in_Dir_HeadVld; // @[router.scala 240:240 242:24 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h2
     : io_Sta_in_Dir_HeadPtr; // @[router.scala 240:240 243:24 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 240:240 244:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_MemData; // @[router.scala 240:240 245:20 node.scala 25:11]
  wire [1:0] _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h1
     : io_Sta_in_HomeProc_CacheState; // @[router.scala 240:240 246:32 node.scala 25:11]
  wire [2:0] _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 3'h3
     : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 240:240 247:28 node.scala 25:11]
  wire [1:0] _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_RpMsg_2_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_UniMsg_2_Data; // @[router.scala 240:240 248:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_5 : io_Sta_in_HomeProc_CacheState; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_0 : io_Sta_in_Dir_Dirty; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadVld; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_en_r ? _GEN_4 : io_Sta_in_MemData; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_6 : io_Sta_in_UniMsg_2_Cmd; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_7 : io_Sta_in_UniMsg_2_Data; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_Get_Put_Dirty_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_Dirty; // @[router.scala 240:240 241:22 node.scala 25:11]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) |
    io_Sta_in_Dir_HeadVld; // @[router.scala 240:240 242:24 node.scala 25:11]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h3
     : io_Sta_in_Dir_HeadPtr; // @[router.scala 240:240 243:24 node.scala 25:11]
  wire  _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 240:240 244:28 node.scala 25:11]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_MemData; // @[router.scala 240:240 245:20 node.scala 25:11]
  wire [1:0] _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 2'h1
     : io_Sta_in_HomeProc_CacheState; // @[router.scala 240:240 246:32 node.scala 25:11]
  wire [2:0] _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ? 3'h3
     : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 240:240 247:28 node.scala 25:11]
  wire [1:0] _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_RpMsg_3_Cmd & (~
    io_Sta_in_Dir_Pending & (io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState == 2'h2))))) ?
    io_Sta_in_HomeProc_CacheData : io_Sta_in_UniMsg_3_Data; // @[router.scala 240:240 248:29 node.scala 25:11]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_5 : io_Sta_in_HomeProc_CacheState; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_0 : io_Sta_in_Dir_Dirty; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_1 : io_Sta_in_Dir_HeadVld; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_en_r ? _GEN_4 : io_Sta_in_MemData; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_6 : io_Sta_in_UniMsg_3_Cmd; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_7 : io_Sta_in_UniMsg_3_Data; // @[router.scala 239:14 node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc &
    io_Sta_in_Proc_2_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc &
    io_Sta_in_Proc_3_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc &
    io_Sta_in_Proc_1_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_4(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc &
    io_Sta_in_Proc_3_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_6(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc &
    io_Sta_in_Proc_1_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_7(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 254:186 255:28]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc &
    io_Sta_in_Proc_2_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 254:186 256:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_8(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 253:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h1 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_1_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 263:27]
  wire  _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h1 & (~io_Sta_in_HomeUniMsg_HomeProc
     & io_Sta_in_Proc_1_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 264:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_0 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_Home_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h2 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_2_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 263:27]
  wire  _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h2 & (~io_Sta_in_HomeUniMsg_HomeProc
     & io_Sta_in_Proc_2_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 264:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_0 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Nak_Home_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h3 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_3_CacheState != 2'h2)) ? 3'h5 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 263:27]
  wire  _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h3 & (~io_Sta_in_HomeUniMsg_HomeProc
     & io_Sta_in_Proc_3_CacheState != 2'h2)) | io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 262:164 264:24]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_0 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11 router.scala 261:14]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? io_Sta_in_Proc_2_CacheData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc &
    io_Sta_in_Proc_2_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h2 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? io_Sta_in_Proc_2_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? io_Sta_in_Proc_3_CacheData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc &
    io_Sta_in_Proc_3_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h1 & (io_Sta_in_UniMsg_1_Proc == 2'h3 & (~io_Sta_in_UniMsg_1_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? io_Sta_in_Proc_3_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? io_Sta_in_Proc_1_CacheData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h2 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc &
    io_Sta_in_Proc_1_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h1 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? io_Sta_in_Proc_1_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_4(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? io_Sta_in_Proc_3_CacheData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h2 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc &
    io_Sta_in_Proc_3_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h1 & (io_Sta_in_UniMsg_2_Proc == 2'h3 & (~io_Sta_in_UniMsg_2_HomeProc
     & io_Sta_in_Proc_3_CacheState == 2'h2)) ? io_Sta_in_Proc_3_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_6(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? io_Sta_in_Proc_1_CacheData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h3 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc &
    io_Sta_in_Proc_1_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h1 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_1_CacheState == 2'h2)) ? io_Sta_in_Proc_1_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_7(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 270:186 271:33]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 270:186 272:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? io_Sta_in_Proc_2_CacheData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 270:186 273:29]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 270:186 274:24]
  wire [1:0] _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h3 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 270:186 275:25]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc &
    io_Sta_in_Proc_2_CacheState == 2'h2)) ? 1'h0 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 270:186 276:29]
  wire [1:0] _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h1 & (io_Sta_in_UniMsg_3_Proc == 2'h2 & (~io_Sta_in_UniMsg_3_HomeProc
     & io_Sta_in_Proc_2_CacheState == 2'h2)) ? io_Sta_in_Proc_2_CacheData : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 270:186 277:25]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_en_r ? _GEN_3 : io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_en_r ? _GEN_4 : io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_en_r ? _GEN_5 : io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_en_r ? _GEN_6 : io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_8(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11 router.scala 269:14]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h1 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 283:164 284:33]
  wire [2:0] _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h1 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_1_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 283:164 285:27]
  wire [1:0] _GEN_2 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h1 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_1_CacheState == 2'h2)) ? io_Sta_in_Proc_1_CacheData :
    io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 283:164 286:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_en_r ? _GEN_2 : io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_Home_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h2 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 283:164 284:33]
  wire [2:0] _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h2 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_2_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 283:164 285:27]
  wire [1:0] _GEN_2 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h2 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_2_CacheState == 2'h2)) ? io_Sta_in_Proc_2_CacheData :
    io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 283:164 286:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_en_r ? _GEN_2 : io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Remote_Get_Put_Home_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [1:0] _GEN_0 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h3 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 2'h1 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 283:164 284:33]
  wire [2:0] _GEN_1 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h3 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_3_CacheState == 2'h2)) ? 3'h3 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 283:164 285:27]
  wire [1:0] _GEN_2 = io_Sta_in_HomeUniMsg_Cmd == 3'h1 & (io_Sta_in_HomeUniMsg_Proc == 2'h3 & (~
    io_Sta_in_HomeUniMsg_HomeProc & io_Sta_in_Proc_3_CacheState == 2'h2)) ? io_Sta_in_Proc_3_CacheData :
    io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 283:164 286:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_en_r ? _GEN_0 : io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_en_r ? _GEN_1 : io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_en_r ? _GEN_2 : io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11 router.scala 282:14]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_Nak(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (io_Sta_in_Dir_Pending | (
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) | io_Sta_in_Dir_Dirty & (~
    io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h1 & ~io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h5 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 292:311 293:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 291:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_Nak_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (io_Sta_in_Dir_Pending | (
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) | io_Sta_in_Dir_Dirty & (~
    io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h2 & ~io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h5 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 292:311 293:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 291:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_Nak_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire [2:0] _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (io_Sta_in_Dir_Pending | (
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_CacheState != 2'h2) | io_Sta_in_Dir_Dirty & (~
    io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr == 2'h3 & ~io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h5 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 292:311 293:28]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_0 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 291:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_GetX(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr))))) |
    io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 299:220 300:24]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h2
     : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 299:220 301:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11 router.scala 299:220 302:29]
  wire  _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 299:220 303:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_1_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_1_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_GetX_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr))))) |
    io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 299:220 300:24]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h2
     : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 299:220 301:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11 router.scala 299:220 302:29]
  wire  _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 299:220 303:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_2_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_2_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_GetX_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr))))) |
    io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 299:220 300:24]
  wire [2:0] _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr))))) ? 3'h2
     : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 299:220 301:28]
  wire [1:0] _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HeadPtr : io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11 router.scala 299:220 302:29]
  wire  _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_Local & (io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr))))) ?
    io_Sta_in_Dir_HomeHeadPtr : io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 299:220 303:33]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_0 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_1 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_3_Proc = io_en_r ? _GEN_2 : io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_3_HomeProc = io_en_r ? _GEN_3 : io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11 router.scala 298:14]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 309:227 310:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 309:227 311:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 309:227 312:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h1
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 309:227 313:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 309:227 314:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 309:227 315:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 309:227 321:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 309:227 322:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 309:227 323:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 309:227 324:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 309:227 325:32]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 309:227 326:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_17 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_1_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 309:227 310:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 309:227 311:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 309:227 312:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h2
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 309:227 313:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 309:227 314:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 309:227 315:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 309:227 321:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 309:227 322:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 309:227 323:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 309:227 324:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 309:227 325:32]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 309:227 326:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_17 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_1_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 309:227 310:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 309:227 311:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 309:227 312:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h3
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 309:227 313:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 309:227 314:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 309:227 315:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 309:227 317:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 309:227 318:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 309:227 321:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 309:227 322:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 309:227 323:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 309:227 324:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 309:227 325:32]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 309:227 326:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_17 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 308:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 332:227 333:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 332:227 334:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 332:227 335:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h1
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 332:227 336:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 332:227 337:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 332:227 338:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 332:227 344:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 332:227 345:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 332:227 346:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 332:227 347:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 332:227 348:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_2_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 332:227 333:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 332:227 334:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 332:227 335:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h2
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 332:227 336:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 332:227 337:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 332:227 338:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 332:227 344:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 332:227 345:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 332:227 346:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 332:227 347:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 332:227 348:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_2_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 332:227 333:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 332:227 334:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) |
    io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 332:227 335:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h3
     : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 332:227 336:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 332:227 337:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 332:227 338:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 332:227 340:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 332:227 341:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 332:227 344:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 1'h0
     : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 332:227 345:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 3'h4
     : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 332:227 346:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ?
    io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 332:227 347:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1))))) ? 2'h0
     : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 332:227 348:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 331:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 354:187 355:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 354:187 356:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 354:187 357:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 354:187 358:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 354:187 359:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 354:187 360:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 354:187 366:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 354:187 367:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 354:187 368:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 354:187 369:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 354:187 370:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_3_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 354:187 355:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 354:187 356:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 354:187 357:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 354:187 358:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 354:187 359:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 354:187 360:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 354:187 366:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 354:187 367:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 354:187 368:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 354:187 369:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 354:187 370:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_3_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _GEN_0 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 354:187 355:22]
  wire  _GEN_1 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 354:187 356:22]
  wire  _GEN_2 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 354:187 357:24]
  wire [1:0] _GEN_3 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 354:187 358:24]
  wire  _GEN_4 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 354:187 359:28]
  wire  _GEN_5 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 354:187 360:23]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 354:187 362:26]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 354:187 363:26]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 354:187 366:27]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 354:187 367:27]
  wire [2:0] _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 3'h4 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 354:187 368:28]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 354:187 369:29]
  wire [1:0] _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (~io_Sta_in_Dir_HeadVld & ~io_Sta_in_Dir_Local)))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 354:187 370:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_16 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_1 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_2 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_4 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_5 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_6 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_8 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_10 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_12 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_7 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_9 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_11 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_13 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_14 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_15 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 353:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_4(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_4_1(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_4_2(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 375:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_5(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_5_1(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_5_2(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 398:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_6(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_6_1(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_6_2(
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_Sta_in_Dir_Pending; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Local = io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_Dirty = io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadVld = io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HeadPtr = io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrVld = io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeShrSet = io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_2 = io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_InvSet_3 = io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_Dir_HomeInvSet = io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 420:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeInvMsg_Cmd = io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_27 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _T_35 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 443:288 444:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 443:288 445:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 443:288 446:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 443:288 447:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 443:288 448:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 443:288 449:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 443:288 450:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_27 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_35 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 443:288 462:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 443:288 463:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 443:288 464:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 443:288 465:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 443:288 466:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 443:288 467:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_19 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _T_35 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 443:288 444:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 443:288 445:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 443:288 446:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 443:288 447:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 443:288 448:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 443:288 449:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 443:288 450:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_19 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_35 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 443:288 462:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 443:288 463:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 443:288 464:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 443:288 465:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 443:288 466:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 443:288 467:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_19 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _T_27 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 453:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 453:161 455:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 443:288 444:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 443:288 445:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 443:288 446:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 443:288 447:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 443:288 448:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 443:288 449:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 443:288 450:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_19 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _T_27 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 443:288]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 443:288 452:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 443:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 443:288 462:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 443:288 463:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 443:288 464:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 443:288 465:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 443:288 466:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 443:288 467:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 442:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7_NODE_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_27 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _T_35 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 473:288 474:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 473:288 475:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 473:288 476:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 473:288 477:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 473:288 478:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 473:288 479:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 473:288 480:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_27 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_35 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 473:288 492:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 473:288 493:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 473:288 494:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 473:288 495:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 473:288 496:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 473:288 497:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 473:288 498:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7_NODE_Get_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_19 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _T_35 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 473:288 474:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 473:288 475:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 473:288 476:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 473:288 477:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 473:288 478:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 473:288 479:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 473:288 480:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_19 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_35 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 473:288 492:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 473:288 493:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 473:288 494:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 473:288 495:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 473:288 496:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 473:288 497:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 473:288 498:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_7_NODE_Get_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_19 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _T_27 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 483:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 483:161 485:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 473:288 474:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 473:288 475:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 473:288 476:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 473:288 477:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 473:288 478:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 473:288 479:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 473:288 480:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_19 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _T_27 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 473:288]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 473:288 482:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 473:288]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 473:288 492:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 473:288 493:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 473:288 494:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 3'h4 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 473:288 495:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 473:288 496:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) ? 2'h0 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 473:288 497:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & (
    io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))) | io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 473:288 498:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 472:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 504:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 504:319 505:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 504:319 506:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 504:319 507:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 504:319 508:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 504:319 509:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 504:319 510:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 504:319 511:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 504:319 523:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 504:319 524:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 504:319 525:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 504:319 526:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 504:319 527:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 504:319 528:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 504:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 504:319 505:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 504:319 506:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 504:319 507:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 504:319 508:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 504:319 509:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 504:319 510:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 504:319 511:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 504:319 523:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 504:319 524:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 504:319 525:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 504:319 526:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 504:319 527:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 504:319 528:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 504:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 514:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 514:161 516:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 504:319 505:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 504:319 506:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 504:319 507:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 504:319 508:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 504:319 509:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 504:319 510:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 504:319 511:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 504:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 504:319 513:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 504:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 504:319 523:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 504:319 524:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 504:319 525:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 504:319 526:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 504:319 527:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 504:319 528:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 503:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home_NODE_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 534:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 534:319 535:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 534:319 536:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 534:319 537:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 534:319 538:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 534:319 539:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 534:319 540:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 534:319 541:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 534:319 553:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 534:319 554:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 534:319 555:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 534:319 556:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 534:319 557:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 534:319 558:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 534:319 559:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home_NODE_Get_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 534:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 534:319 535:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 534:319 536:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 534:319 537:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 534:319 538:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 534:319 539:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 534:319 540:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 534:319 541:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 534:319 553:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 534:319 554:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 534:319 555:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 534:319 556:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 534:319 557:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 534:319 558:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 534:319 559:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_Home_NODE_Get_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 534:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 544:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 544:161 546:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending
    ; // @[node.scala 25:11 router.scala 534:319 535:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 534:319 536:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 534:319 537:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld
    ; // @[node.scala 25:11 router.scala 534:319 538:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 534:319 539:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 534:319 540:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 534:319 541:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 534:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 534:319 543:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 534:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 534:319 553:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 534:319 554:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 534:319 555:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 534:319 556:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 534:319 557:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 534:319 558:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 534:319 559:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 533:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_4(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_6(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_7(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_8(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 565:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 575:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 575:161 577:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 565:319 566:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 565:319 567:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 565:319 568:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 565:319 569:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 565:319 570:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 565:319 571:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 565:319 572:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 565:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 565:319 574:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 565:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 565:319 584:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 565:319 585:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 565:319 586:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 565:319 587:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 565:319 588:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd != 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 565:319 589:32]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 564:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h1 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_4(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_37 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h2 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_37 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_5 :
    io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_6(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_7(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_8_NODE_Get_8(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 595:192]
  wire  _T_21 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _T_29 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 605:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 605:161 607:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 595:319 596:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 595:319 597:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 595:319 598:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 595:319 599:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h3 :
    io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 595:319 600:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 595:319 601:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 595:319 602:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_21 :
    io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_1 :
    io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _T_29 :
    io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 595:319]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? _GEN_3 :
    io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 595:319 604:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 595:319]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 595:319 614:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 1'h0 :
    io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 595:319 615:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 595:319 616:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 3'h4 :
    io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 595:319 617:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? io_Sta_in_MemData :
    io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 595:319 618:29]
  wire [1:0] _GEN_27 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) ? 2'h0 :
    io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 595:319 619:32]
  wire  _GEN_28 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & (io_Sta_in_Dir_Local & io_Sta_in_HomeProc_ProcCmd == 2'h1)))))))) |
    io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 595:319 620:31]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_en_r ? _GEN_28 : io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheState = io_en_r ? _GEN_27 : io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 594:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_9(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_26 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _T_34 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 626:248 627:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 626:248 628:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 626:248 629:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 626:248 630:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 626:248 631:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 626:248 632:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 626:248 633:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_26 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_34 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 626:248 645:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 626:248 646:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 626:248 647:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 626:248 648:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h1 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 626:248 649:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_9_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_18 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _T_34 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 626:248 627:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 626:248 628:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 626:248 629:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 626:248 630:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 626:248 631:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 626:248 632:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 626:248 633:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_18 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_34 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 626:248 645:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 626:248 646:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 626:248 647:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 626:248 648:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h2 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 626:248 649:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_9_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_18 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _T_26 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr); // @[router.scala 636:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & ~io_Sta_in_Dir_HomeHeadPtr) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 636:161 638:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 626:248 627:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 626:248 628:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 626:248 629:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 626:248 630:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 626:248 631:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 626:248 632:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 626:248 633:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_18 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _T_26 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 626:248]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 626:248 635:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 626:248]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 626:248 645:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 626:248 646:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 626:248 647:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? 3'h4 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 626:248 648:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & ((io_Sta_in_Dir_HeadPtr != 2'h3 | io_Sta_in_Dir_HomeHeadPtr) & ~
    io_Sta_in_Dir_Local))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 626:248 649:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 625:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_Home(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 655:192]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 655:279 656:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 655:279 657:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 655:279 658:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 655:279 659:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 655:279 660:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 655:279 661:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 655:279 662:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 655:279 674:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 655:279 675:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 655:279 676:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 655:279 677:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 655:279 678:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_Home_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 655:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 655:279 656:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 655:279 657:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 655:279 658:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 655:279 659:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 655:279 660:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 655:279 661:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 655:279 662:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 655:279 674:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 655:279 675:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 655:279 676:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 655:279 677:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 655:279 678:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_Home_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 655:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 665:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 665:161 667:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 655:279 656:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 655:279 657:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 655:279 658:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 655:279 659:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 655:279 660:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 655:279 661:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 655:279 662:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 655:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 655:279 664:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 655:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 655:279 674:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 655:279 675:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 655:279 676:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 655:279 677:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_HomeShrSet & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 655:279 678:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 654:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_1(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_2(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 2'h1 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_1_Cmd == 3'h2 & (io_Sta_in_UniMsg_1_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Cmd = io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_en_r ? _GEN_18 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_3(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_4(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_2 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_5(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_36 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_5 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_3 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 2'h2 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _T_36 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_21 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? _GEN_5 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_22 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 684:279 703:27]
  wire  _GEN_23 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 684:279 704:27]
  wire [1:0] _GEN_24 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 2'h0 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 684:279 705:27]
  wire [2:0] _GEN_25 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? 3'h4 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279 706:28]
  wire [1:0] _GEN_26 = io_Sta_in_UniMsg_2_Cmd == 3'h2 & (io_Sta_in_UniMsg_2_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_3 & ~io_Sta_in_Dir_Local))))))) ? io_Sta_in_MemData : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 684:279 707:29]
  assign io_Sta_out_Proc_0_ProcCmd = io_Sta_in_Proc_0_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_InvMarked = io_Sta_in_Proc_0_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheState = io_Sta_in_Proc_0_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_0_CacheData = io_Sta_in_Proc_0_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_ProcCmd = io_Sta_in_Proc_1_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_InvMarked = io_Sta_in_Proc_1_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheState = io_Sta_in_Proc_1_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_1_CacheData = io_Sta_in_Proc_1_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_ProcCmd = io_Sta_in_Proc_2_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_InvMarked = io_Sta_in_Proc_2_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheState = io_Sta_in_Proc_2_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_2_CacheData = io_Sta_in_Proc_2_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_ProcCmd = io_Sta_in_Proc_3_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_InvMarked = io_Sta_in_Proc_3_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheState = io_Sta_in_Proc_3_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_Proc_3_CacheData = io_Sta_in_Proc_3_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_ProcCmd = io_Sta_in_HomeProc_ProcCmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_InvMarked = io_Sta_in_HomeProc_InvMarked; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheState = io_Sta_in_HomeProc_CacheState; // @[node.scala 25:11]
  assign io_Sta_out_HomeProc_CacheData = io_Sta_in_HomeProc_CacheData; // @[node.scala 25:11]
  assign io_Sta_out_Dir_Pending = io_en_r ? _GEN_6 : io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Local = io_en_r ? _GEN_7 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_Dirty = io_en_r ? _GEN_8 : io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadVld = io_en_r ? _GEN_9 : io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HeadPtr = io_en_r ? _GEN_10 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeHeadPtr = io_en_r ? _GEN_11 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrVld = io_en_r ? _GEN_12 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_0 = io_Sta_in_Dir_ShrSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_ShrSet_1 = io_en_r ? _GEN_13 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_2 = io_en_r ? _GEN_16 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_ShrSet_3 = io_en_r ? _GEN_19 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeShrSet = io_en_r ? _GEN_22 : io_Sta_in_Dir_HomeShrSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_0 = io_Sta_in_Dir_InvSet_0; // @[node.scala 25:11]
  assign io_Sta_out_Dir_InvSet_1 = io_en_r ? _GEN_14 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_2 = io_en_r ? _GEN_17 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_InvSet_3 = io_en_r ? _GEN_20 : io_Sta_in_Dir_InvSet_3; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_Dir_HomeInvSet = io_en_r ? _GEN_23 : io_Sta_in_Dir_HomeInvSet; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_MemData = io_Sta_in_MemData; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Cmd = io_Sta_in_UniMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Proc = io_Sta_in_UniMsg_0_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_HomeProc = io_Sta_in_UniMsg_0_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_0_Data = io_Sta_in_UniMsg_0_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Cmd = io_Sta_in_UniMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Proc = io_Sta_in_UniMsg_1_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_HomeProc = io_Sta_in_UniMsg_1_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_1_Data = io_Sta_in_UniMsg_1_Data; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Cmd = io_en_r ? _GEN_25 : io_Sta_in_UniMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_2_Proc = io_Sta_in_UniMsg_2_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_HomeProc = io_Sta_in_UniMsg_2_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_2_Data = io_en_r ? _GEN_26 : io_Sta_in_UniMsg_2_Data; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_UniMsg_3_Cmd = io_Sta_in_UniMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Proc = io_Sta_in_UniMsg_3_Proc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_HomeProc = io_Sta_in_UniMsg_3_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_UniMsg_3_Data = io_Sta_in_UniMsg_3_Data; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Cmd = io_Sta_in_HomeUniMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Proc = io_Sta_in_HomeUniMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_HomeProc = io_Sta_in_HomeUniMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_HomeUniMsg_Data = io_Sta_in_HomeUniMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_0_Cmd = io_Sta_in_InvMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_InvMsg_1_Cmd = io_en_r ? _GEN_15 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_2_Cmd = io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_InvMsg_3_Cmd = io_en_r ? _GEN_21 : io_Sta_in_InvMsg_3_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_HomeInvMsg_Cmd = io_en_r ? _GEN_24 : io_Sta_in_HomeInvMsg_Cmd; // @[node.scala 25:11 router.scala 683:14]
  assign io_Sta_out_RpMsg_0_Cmd = io_Sta_in_RpMsg_0_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_1_Cmd = io_Sta_in_RpMsg_1_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_2_Cmd = io_Sta_in_RpMsg_2_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_RpMsg_3_Cmd = io_Sta_in_RpMsg_3_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_HomeRpMsg_Cmd = io_Sta_in_HomeRpMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Cmd = io_Sta_in_WbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Proc = io_Sta_in_WbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_HomeProc = io_Sta_in_WbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_WbMsg_Data = io_Sta_in_WbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Cmd = io_Sta_in_ShWbMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Proc = io_Sta_in_ShWbMsg_Proc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_HomeProc = io_Sta_in_ShWbMsg_HomeProc; // @[node.scala 25:11]
  assign io_Sta_out_ShWbMsg_Data = io_Sta_in_ShWbMsg_Data; // @[node.scala 25:11]
  assign io_Sta_out_NakcMsg_Cmd = io_Sta_in_NakcMsg_Cmd; // @[node.scala 25:11]
  assign io_Sta_out_CurrData = io_Sta_in_CurrData; // @[node.scala 25:11]
endmodule
module NI_Local_GetX_PutX_10_6(
  input        io_en_r,
  input  [1:0] io_Sta_in_Proc_0_ProcCmd,
  input        io_Sta_in_Proc_0_InvMarked,
  input  [1:0] io_Sta_in_Proc_0_CacheState,
  input  [1:0] io_Sta_in_Proc_0_CacheData,
  input  [1:0] io_Sta_in_Proc_1_ProcCmd,
  input        io_Sta_in_Proc_1_InvMarked,
  input  [1:0] io_Sta_in_Proc_1_CacheState,
  input  [1:0] io_Sta_in_Proc_1_CacheData,
  input  [1:0] io_Sta_in_Proc_2_ProcCmd,
  input        io_Sta_in_Proc_2_InvMarked,
  input  [1:0] io_Sta_in_Proc_2_CacheState,
  input  [1:0] io_Sta_in_Proc_2_CacheData,
  input  [1:0] io_Sta_in_Proc_3_ProcCmd,
  input        io_Sta_in_Proc_3_InvMarked,
  input  [1:0] io_Sta_in_Proc_3_CacheState,
  input  [1:0] io_Sta_in_Proc_3_CacheData,
  input  [1:0] io_Sta_in_HomeProc_ProcCmd,
  input        io_Sta_in_HomeProc_InvMarked,
  input  [1:0] io_Sta_in_HomeProc_CacheState,
  input  [1:0] io_Sta_in_HomeProc_CacheData,
  input        io_Sta_in_Dir_Pending,
  input        io_Sta_in_Dir_Local,
  input        io_Sta_in_Dir_Dirty,
  input        io_Sta_in_Dir_HeadVld,
  input  [1:0] io_Sta_in_Dir_HeadPtr,
  input        io_Sta_in_Dir_HomeHeadPtr,
  input        io_Sta_in_Dir_ShrVld,
  input        io_Sta_in_Dir_ShrSet_0,
  input        io_Sta_in_Dir_ShrSet_1,
  input        io_Sta_in_Dir_ShrSet_2,
  input        io_Sta_in_Dir_ShrSet_3,
  input        io_Sta_in_Dir_HomeShrSet,
  input        io_Sta_in_Dir_InvSet_0,
  input        io_Sta_in_Dir_InvSet_1,
  input        io_Sta_in_Dir_InvSet_2,
  input        io_Sta_in_Dir_InvSet_3,
  input        io_Sta_in_Dir_HomeInvSet,
  input  [1:0] io_Sta_in_MemData,
  input  [2:0] io_Sta_in_UniMsg_0_Cmd,
  input  [1:0] io_Sta_in_UniMsg_0_Proc,
  input        io_Sta_in_UniMsg_0_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_0_Data,
  input  [2:0] io_Sta_in_UniMsg_1_Cmd,
  input  [1:0] io_Sta_in_UniMsg_1_Proc,
  input        io_Sta_in_UniMsg_1_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_1_Data,
  input  [2:0] io_Sta_in_UniMsg_2_Cmd,
  input  [1:0] io_Sta_in_UniMsg_2_Proc,
  input        io_Sta_in_UniMsg_2_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_2_Data,
  input  [2:0] io_Sta_in_UniMsg_3_Cmd,
  input  [1:0] io_Sta_in_UniMsg_3_Proc,
  input        io_Sta_in_UniMsg_3_HomeProc,
  input  [1:0] io_Sta_in_UniMsg_3_Data,
  input  [2:0] io_Sta_in_HomeUniMsg_Cmd,
  input  [1:0] io_Sta_in_HomeUniMsg_Proc,
  input        io_Sta_in_HomeUniMsg_HomeProc,
  input  [1:0] io_Sta_in_HomeUniMsg_Data,
  input  [1:0] io_Sta_in_InvMsg_0_Cmd,
  input  [1:0] io_Sta_in_InvMsg_1_Cmd,
  input  [1:0] io_Sta_in_InvMsg_2_Cmd,
  input  [1:0] io_Sta_in_InvMsg_3_Cmd,
  input  [1:0] io_Sta_in_HomeInvMsg_Cmd,
  input        io_Sta_in_RpMsg_0_Cmd,
  input        io_Sta_in_RpMsg_1_Cmd,
  input        io_Sta_in_RpMsg_2_Cmd,
  input        io_Sta_in_RpMsg_3_Cmd,
  input        io_Sta_in_HomeRpMsg_Cmd,
  input        io_Sta_in_WbMsg_Cmd,
  input  [1:0] io_Sta_in_WbMsg_Proc,
  input        io_Sta_in_WbMsg_HomeProc,
  input  [1:0] io_Sta_in_WbMsg_Data,
  input  [1:0] io_Sta_in_ShWbMsg_Cmd,
  input  [1:0] io_Sta_in_ShWbMsg_Proc,
  input        io_Sta_in_ShWbMsg_HomeProc,
  input  [1:0] io_Sta_in_ShWbMsg_Data,
  input        io_Sta_in_NakcMsg_Cmd,
  input  [1:0] io_Sta_in_CurrData,
  output [1:0] io_Sta_out_Proc_0_ProcCmd,
  output       io_Sta_out_Proc_0_InvMarked,
  output [1:0] io_Sta_out_Proc_0_CacheState,
  output [1:0] io_Sta_out_Proc_0_CacheData,
  output [1:0] io_Sta_out_Proc_1_ProcCmd,
  output       io_Sta_out_Proc_1_InvMarked,
  output [1:0] io_Sta_out_Proc_1_CacheState,
  output [1:0] io_Sta_out_Proc_1_CacheData,
  output [1:0] io_Sta_out_Proc_2_ProcCmd,
  output       io_Sta_out_Proc_2_InvMarked,
  output [1:0] io_Sta_out_Proc_2_CacheState,
  output [1:0] io_Sta_out_Proc_2_CacheData,
  output [1:0] io_Sta_out_Proc_3_ProcCmd,
  output       io_Sta_out_Proc_3_InvMarked,
  output [1:0] io_Sta_out_Proc_3_CacheState,
  output [1:0] io_Sta_out_Proc_3_CacheData,
  output [1:0] io_Sta_out_HomeProc_ProcCmd,
  output       io_Sta_out_HomeProc_InvMarked,
  output [1:0] io_Sta_out_HomeProc_CacheState,
  output [1:0] io_Sta_out_HomeProc_CacheData,
  output       io_Sta_out_Dir_Pending,
  output       io_Sta_out_Dir_Local,
  output       io_Sta_out_Dir_Dirty,
  output       io_Sta_out_Dir_HeadVld,
  output [1:0] io_Sta_out_Dir_HeadPtr,
  output       io_Sta_out_Dir_HomeHeadPtr,
  output       io_Sta_out_Dir_ShrVld,
  output       io_Sta_out_Dir_ShrSet_0,
  output       io_Sta_out_Dir_ShrSet_1,
  output       io_Sta_out_Dir_ShrSet_2,
  output       io_Sta_out_Dir_ShrSet_3,
  output       io_Sta_out_Dir_HomeShrSet,
  output       io_Sta_out_Dir_InvSet_0,
  output       io_Sta_out_Dir_InvSet_1,
  output       io_Sta_out_Dir_InvSet_2,
  output       io_Sta_out_Dir_InvSet_3,
  output       io_Sta_out_Dir_HomeInvSet,
  output [1:0] io_Sta_out_MemData,
  output [2:0] io_Sta_out_UniMsg_0_Cmd,
  output [1:0] io_Sta_out_UniMsg_0_Proc,
  output       io_Sta_out_UniMsg_0_HomeProc,
  output [1:0] io_Sta_out_UniMsg_0_Data,
  output [2:0] io_Sta_out_UniMsg_1_Cmd,
  output [1:0] io_Sta_out_UniMsg_1_Proc,
  output       io_Sta_out_UniMsg_1_HomeProc,
  output [1:0] io_Sta_out_UniMsg_1_Data,
  output [2:0] io_Sta_out_UniMsg_2_Cmd,
  output [1:0] io_Sta_out_UniMsg_2_Proc,
  output       io_Sta_out_UniMsg_2_HomeProc,
  output [1:0] io_Sta_out_UniMsg_2_Data,
  output [2:0] io_Sta_out_UniMsg_3_Cmd,
  output [1:0] io_Sta_out_UniMsg_3_Proc,
  output       io_Sta_out_UniMsg_3_HomeProc,
  output [1:0] io_Sta_out_UniMsg_3_Data,
  output [2:0] io_Sta_out_HomeUniMsg_Cmd,
  output [1:0] io_Sta_out_HomeUniMsg_Proc,
  output       io_Sta_out_HomeUniMsg_HomeProc,
  output [1:0] io_Sta_out_HomeUniMsg_Data,
  output [1:0] io_Sta_out_InvMsg_0_Cmd,
  output [1:0] io_Sta_out_InvMsg_1_Cmd,
  output [1:0] io_Sta_out_InvMsg_2_Cmd,
  output [1:0] io_Sta_out_InvMsg_3_Cmd,
  output [1:0] io_Sta_out_HomeInvMsg_Cmd,
  output       io_Sta_out_RpMsg_0_Cmd,
  output       io_Sta_out_RpMsg_1_Cmd,
  output       io_Sta_out_RpMsg_2_Cmd,
  output       io_Sta_out_RpMsg_3_Cmd,
  output       io_Sta_out_HomeRpMsg_Cmd,
  output       io_Sta_out_WbMsg_Cmd,
  output [1:0] io_Sta_out_WbMsg_Proc,
  output       io_Sta_out_WbMsg_HomeProc,
  output [1:0] io_Sta_out_WbMsg_Data,
  output [1:0] io_Sta_out_ShWbMsg_Cmd,
  output [1:0] io_Sta_out_ShWbMsg_Proc,
  output       io_Sta_out_ShWbMsg_HomeProc,
  output [1:0] io_Sta_out_ShWbMsg_Data,
  output       io_Sta_out_NakcMsg_Cmd,
  output [1:0] io_Sta_out_CurrData
);
  wire  _T_4 = ~io_Sta_in_Dir_HomeHeadPtr; // @[router.scala 684:192]
  wire  _T_20 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_1 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_1 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h1
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _T_28 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4); // @[router.scala 694:70]
  wire [1:0] _GEN_3 = io_Sta_in_Dir_ShrVld & io_Sta_in_Dir_ShrSet_2 | io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h2
     & _T_4) ? 2'h1 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 694:161 696:26]
  wire  _GEN_6 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Pending; // @[node.scala 25:11 router.scala 684:279 685:24]
  wire  _GEN_7 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_Local; // @[node.scala 25:11 router.scala 684:279 686:22]
  wire  _GEN_8 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_Dirty; // @[node.scala 25:11 router.scala 684:279 687:22]
  wire  _GEN_9 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) | io_Sta_in_Dir_HeadVld; // @[node.scala 25:11 router.scala 684:279 688:24]
  wire [1:0] _GEN_10 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 2'h3 : io_Sta_in_Dir_HeadPtr; // @[node.scala 25:11 router.scala 684:279 689:24]
  wire  _GEN_11 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_HomeHeadPtr; // @[node.scala 25:11 router.scala 684:279 690:28]
  wire  _GEN_12 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrVld; // @[node.scala 25:11 router.scala 684:279 691:23]
  wire  _GEN_13 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_1; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_14 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_20 : io_Sta_in_Dir_InvSet_1; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_15 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_1 : io_Sta_in_InvMsg_1_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_16 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_2; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_17 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _T_28 : io_Sta_in_Dir_InvSet_2; // @[node.scala 25:11 router.scala 684:279]
  wire [1:0] _GEN_18 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? _GEN_3 : io_Sta_in_InvMsg_2_Cmd; // @[node.scala 25:11 router.scala 684:279]
  wire  _GEN_19 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
    io_Sta_in_Dir_ShrSet_1 & ~io_Sta_in_Dir_Local))))))) ? 1'h0 : io_Sta_in_Dir_ShrSet_3; // @[node.scala 25:11 router.scala 684:279 693:26]
  wire  _GEN_20 = io_Sta_in_UniMsg_3_Cmd == 3'h2 & (io_Sta_in_UniMsg_3_HomeProc & (~io_Sta_in_Dir_Pending & (~
    io_Sta_in_Dir_Dirty & (io_Sta_in_Dir_HeadVld & (io_Sta_in_Dir_HeadPtr == 2'h3 & (~io_Sta_in_Dir_HomeHeadPtr & (
