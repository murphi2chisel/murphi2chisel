module Try(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nI_in_1 ? 1'h0 : io_nI_in_1; // @[node.scala 26:10 router.scala 5:18 6:14]
  wire  _GEN_1 = io_nI_in_1 | io_nT_in_1; // @[node.scala 27:10 router.scala 5:18 7:14]
  assign io_x_out = io_x_in; // @[node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_en_r ? _GEN_0 : io_nI_in_1; // @[node.scala 26:10 router.scala 4:14]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_en_r ? _GEN_1 : io_nT_in_1; // @[node.scala 27:10 router.scala 4:14]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Try_1(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nI_in_2 ? 1'h0 : io_nI_in_2; // @[node.scala 26:10 router.scala 5:18 6:14]
  wire  _GEN_1 = io_nI_in_2 | io_nT_in_2; // @[node.scala 27:10 router.scala 5:18 7:14]
  assign io_x_out = io_x_in; // @[node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_en_r ? _GEN_0 : io_nI_in_2; // @[node.scala 26:10 router.scala 4:14]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_en_r ? _GEN_1 : io_nT_in_2; // @[node.scala 27:10 router.scala 4:14]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Crit(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nT_in_1 & io_x_in ? 1'h0 : io_nT_in_1; // @[router.scala 13:40 14:14 node.scala 27:10]
  wire  _GEN_1 = io_nT_in_1 & io_x_in | io_nC_in_1; // @[router.scala 13:40 15:14 node.scala 28:10]
  wire  _GEN_2 = io_nT_in_1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 13:40 16:10 node.scala 25:9]
  assign io_x_out = io_en_r ? _GEN_2 : io_x_in; // @[router.scala 12:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_en_r ? _GEN_0 : io_nT_in_1; // @[router.scala 12:14 node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_en_r ? _GEN_1 : io_nC_in_1; // @[router.scala 12:14 node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Crit_1(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nT_in_2 & io_x_in ? 1'h0 : io_nT_in_2; // @[router.scala 13:40 14:14 node.scala 27:10]
  wire  _GEN_1 = io_nT_in_2 & io_x_in | io_nC_in_2; // @[router.scala 13:40 15:14 node.scala 28:10]
  wire  _GEN_2 = io_nT_in_2 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 13:40 16:10 node.scala 25:9]
  assign io_x_out = io_en_r ? _GEN_2 : io_x_in; // @[router.scala 12:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_en_r ? _GEN_0 : io_nT_in_2; // @[router.scala 12:14 node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_en_r ? _GEN_1 : io_nC_in_2; // @[router.scala 12:14 node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Exit(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nC_in_1 ? 1'h0 : io_nC_in_1; // @[router.scala 22:18 23:14 node.scala 28:10]
  wire  _GEN_1 = io_nC_in_1 | io_nE_in_1; // @[router.scala 22:18 24:14 node.scala 29:10]
  assign io_x_out = io_x_in; // @[node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_en_r ? _GEN_0 : io_nC_in_1; // @[router.scala 21:14 node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_en_r ? _GEN_1 : io_nE_in_1; // @[router.scala 21:14 node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Exit_1(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nC_in_2 ? 1'h0 : io_nC_in_2; // @[router.scala 22:18 23:14 node.scala 28:10]
  wire  _GEN_1 = io_nC_in_2 | io_nE_in_2; // @[router.scala 22:18 24:14 node.scala 29:10]
  assign io_x_out = io_x_in; // @[node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_en_r ? _GEN_0 : io_nC_in_2; // @[router.scala 21:14 node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_en_r ? _GEN_1 : io_nE_in_2; // @[router.scala 21:14 node.scala 29:10]
endmodule
module Idle(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nE_in_1 ? 1'h0 : io_nE_in_1; // @[node.scala 29:10 router.scala 30:18 31:14]
  wire  _GEN_1 = io_nE_in_1 | io_nI_in_1; // @[node.scala 26:10 router.scala 30:18 32:14]
  wire  _GEN_2 = io_nE_in_1 | io_x_in; // @[router.scala 30:18 33:10 node.scala 25:9]
  assign io_x_out = io_en_r ? _GEN_2 : io_x_in; // @[router.scala 29:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_en_r ? _GEN_1 : io_nI_in_1; // @[node.scala 26:10 router.scala 29:14]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_en_r ? _GEN_0 : io_nE_in_1; // @[node.scala 29:10 router.scala 29:14]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Idle_1(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_nE_in_2 ? 1'h0 : io_nE_in_2; // @[node.scala 29:10 router.scala 30:18 31:14]
  wire  _GEN_1 = io_nE_in_2 | io_nI_in_2; // @[node.scala 26:10 router.scala 30:18 32:14]
  wire  _GEN_2 = io_nE_in_2 | io_x_in; // @[router.scala 30:18 33:10 node.scala 25:9]
  assign io_x_out = io_en_r ? _GEN_2 : io_x_in; // @[router.scala 29:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_en_r ? _GEN_1 : io_nI_in_2; // @[node.scala 26:10 router.scala 29:14]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_en_r ? _GEN_0 : io_nE_in_2; // @[node.scala 29:10 router.scala 29:14]
endmodule
module Str_Idle(
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  assign io_x_out = io_x_in; // @[router.scala 38:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module Str_Crit(
  input   io_en_r,
  input   io_x_in,
  output  io_x_out,
  input   io_nI_in_0,
  input   io_nI_in_1,
  input   io_nI_in_2,
  output  io_nI_out_0,
  output  io_nI_out_1,
  output  io_nI_out_2,
  input   io_nT_in_0,
  input   io_nT_in_1,
  input   io_nT_in_2,
  output  io_nT_out_0,
  output  io_nT_out_1,
  output  io_nT_out_2,
  input   io_nC_in_0,
  input   io_nC_in_1,
  input   io_nC_in_2,
  output  io_nC_out_0,
  output  io_nC_out_1,
  output  io_nC_out_2,
  input   io_nE_in_0,
  input   io_nE_in_1,
  input   io_nE_in_2,
  output  io_nE_out_0,
  output  io_nE_out_1,
  output  io_nE_out_2
);
  wire  _GEN_0 = io_x_in ? 1'h0 : io_x_in; // @[router.scala 46:25 47:10 node.scala 25:9]
  assign io_x_out = io_en_r ? _GEN_0 : io_x_in; // @[router.scala 45:14 node.scala 25:9]
  assign io_nI_out_0 = io_nI_in_0; // @[node.scala 26:10]
  assign io_nI_out_1 = io_nI_in_1; // @[node.scala 26:10]
  assign io_nI_out_2 = io_nI_in_2; // @[node.scala 26:10]
  assign io_nT_out_0 = io_nT_in_0; // @[node.scala 27:10]
  assign io_nT_out_1 = io_nT_in_1; // @[node.scala 27:10]
  assign io_nT_out_2 = io_nT_in_2; // @[node.scala 27:10]
  assign io_nC_out_0 = io_nC_in_0; // @[node.scala 28:10]
  assign io_nC_out_1 = io_nC_in_1; // @[node.scala 28:10]
  assign io_nC_out_2 = io_nC_in_2; // @[node.scala 28:10]
  assign io_nE_out_0 = io_nE_in_0; // @[node.scala 29:10]
  assign io_nE_out_1 = io_nE_in_1; // @[node.scala 29:10]
  assign io_nE_out_2 = io_nE_in_2; // @[node.scala 29:10]
endmodule
module system(
  input        clock,
  input        reset,
  input  [3:0] io_en_a,
  output       io_x_out,
  output       io_nI_out_0,
  output       io_nI_out_1,
  output       io_nI_out_2,
  output       io_nT_out_0,
  output       io_nT_out_1,
  output       io_nT_out_2,
  output       io_nC_out_0,
  output       io_nC_out_1,
  output       io_nC_out_2,
  output       io_nE_out_0,
  output       io_nE_out_1,
  output       io_nE_out_2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  rules_0_io_en_r; // @[system.scala 37:16]
  wire  rules_0_io_x_in; // @[system.scala 37:16]
  wire  rules_0_io_x_out; // @[system.scala 37:16]
  wire  rules_0_io_nI_in_0; // @[system.scala 37:16]
  wire  rules_0_io_nI_in_1; // @[system.scala 37:16]
  wire  rules_0_io_nI_in_2; // @[system.scala 37:16]
  wire  rules_0_io_nI_out_0; // @[system.scala 37:16]
  wire  rules_0_io_nI_out_1; // @[system.scala 37:16]
  wire  rules_0_io_nI_out_2; // @[system.scala 37:16]
  wire  rules_0_io_nT_in_0; // @[system.scala 37:16]
  wire  rules_0_io_nT_in_1; // @[system.scala 37:16]
  wire  rules_0_io_nT_in_2; // @[system.scala 37:16]
  wire  rules_0_io_nT_out_0; // @[system.scala 37:16]
  wire  rules_0_io_nT_out_1; // @[system.scala 37:16]
  wire  rules_0_io_nT_out_2; // @[system.scala 37:16]
  wire  rules_0_io_nC_in_0; // @[system.scala 37:16]
  wire  rules_0_io_nC_in_1; // @[system.scala 37:16]
  wire  rules_0_io_nC_in_2; // @[system.scala 37:16]
  wire  rules_0_io_nC_out_0; // @[system.scala 37:16]
  wire  rules_0_io_nC_out_1; // @[system.scala 37:16]
  wire  rules_0_io_nC_out_2; // @[system.scala 37:16]
  wire  rules_0_io_nE_in_0; // @[system.scala 37:16]
  wire  rules_0_io_nE_in_1; // @[system.scala 37:16]
  wire  rules_0_io_nE_in_2; // @[system.scala 37:16]
  wire  rules_0_io_nE_out_0; // @[system.scala 37:16]
  wire  rules_0_io_nE_out_1; // @[system.scala 37:16]
  wire  rules_0_io_nE_out_2; // @[system.scala 37:16]
  wire  rules_1_io_en_r; // @[system.scala 37:16]
  wire  rules_1_io_x_in; // @[system.scala 37:16]
  wire  rules_1_io_x_out; // @[system.scala 37:16]
  wire  rules_1_io_nI_in_0; // @[system.scala 37:16]
  wire  rules_1_io_nI_in_1; // @[system.scala 37:16]
  wire  rules_1_io_nI_in_2; // @[system.scala 37:16]
  wire  rules_1_io_nI_out_0; // @[system.scala 37:16]
  wire  rules_1_io_nI_out_1; // @[system.scala 37:16]
  wire  rules_1_io_nI_out_2; // @[system.scala 37:16]
  wire  rules_1_io_nT_in_0; // @[system.scala 37:16]
  wire  rules_1_io_nT_in_1; // @[system.scala 37:16]
  wire  rules_1_io_nT_in_2; // @[system.scala 37:16]
  wire  rules_1_io_nT_out_0; // @[system.scala 37:16]
  wire  rules_1_io_nT_out_1; // @[system.scala 37:16]
  wire  rules_1_io_nT_out_2; // @[system.scala 37:16]
  wire  rules_1_io_nC_in_0; // @[system.scala 37:16]
  wire  rules_1_io_nC_in_1; // @[system.scala 37:16]
  wire  rules_1_io_nC_in_2; // @[system.scala 37:16]
  wire  rules_1_io_nC_out_0; // @[system.scala 37:16]
  wire  rules_1_io_nC_out_1; // @[system.scala 37:16]
  wire  rules_1_io_nC_out_2; // @[system.scala 37:16]
  wire  rules_1_io_nE_in_0; // @[system.scala 37:16]
  wire  rules_1_io_nE_in_1; // @[system.scala 37:16]
  wire  rules_1_io_nE_in_2; // @[system.scala 37:16]
  wire  rules_1_io_nE_out_0; // @[system.scala 37:16]
  wire  rules_1_io_nE_out_1; // @[system.scala 37:16]
  wire  rules_1_io_nE_out_2; // @[system.scala 37:16]
  wire  rules_2_io_en_r; // @[system.scala 40:16]
  wire  rules_2_io_x_in; // @[system.scala 40:16]
  wire  rules_2_io_x_out; // @[system.scala 40:16]
  wire  rules_2_io_nI_in_0; // @[system.scala 40:16]
  wire  rules_2_io_nI_in_1; // @[system.scala 40:16]
  wire  rules_2_io_nI_in_2; // @[system.scala 40:16]
  wire  rules_2_io_nI_out_0; // @[system.scala 40:16]
  wire  rules_2_io_nI_out_1; // @[system.scala 40:16]
  wire  rules_2_io_nI_out_2; // @[system.scala 40:16]
  wire  rules_2_io_nT_in_0; // @[system.scala 40:16]
  wire  rules_2_io_nT_in_1; // @[system.scala 40:16]
  wire  rules_2_io_nT_in_2; // @[system.scala 40:16]
  wire  rules_2_io_nT_out_0; // @[system.scala 40:16]
  wire  rules_2_io_nT_out_1; // @[system.scala 40:16]
  wire  rules_2_io_nT_out_2; // @[system.scala 40:16]
  wire  rules_2_io_nC_in_0; // @[system.scala 40:16]
  wire  rules_2_io_nC_in_1; // @[system.scala 40:16]
  wire  rules_2_io_nC_in_2; // @[system.scala 40:16]
  wire  rules_2_io_nC_out_0; // @[system.scala 40:16]
  wire  rules_2_io_nC_out_1; // @[system.scala 40:16]
  wire  rules_2_io_nC_out_2; // @[system.scala 40:16]
  wire  rules_2_io_nE_in_0; // @[system.scala 40:16]
  wire  rules_2_io_nE_in_1; // @[system.scala 40:16]
  wire  rules_2_io_nE_in_2; // @[system.scala 40:16]
  wire  rules_2_io_nE_out_0; // @[system.scala 40:16]
  wire  rules_2_io_nE_out_1; // @[system.scala 40:16]
  wire  rules_2_io_nE_out_2; // @[system.scala 40:16]
  wire  rules_3_io_en_r; // @[system.scala 40:16]
  wire  rules_3_io_x_in; // @[system.scala 40:16]
  wire  rules_3_io_x_out; // @[system.scala 40:16]
  wire  rules_3_io_nI_in_0; // @[system.scala 40:16]
  wire  rules_3_io_nI_in_1; // @[system.scala 40:16]
  wire  rules_3_io_nI_in_2; // @[system.scala 40:16]
  wire  rules_3_io_nI_out_0; // @[system.scala 40:16]
  wire  rules_3_io_nI_out_1; // @[system.scala 40:16]
  wire  rules_3_io_nI_out_2; // @[system.scala 40:16]
  wire  rules_3_io_nT_in_0; // @[system.scala 40:16]
  wire  rules_3_io_nT_in_1; // @[system.scala 40:16]
  wire  rules_3_io_nT_in_2; // @[system.scala 40:16]
  wire  rules_3_io_nT_out_0; // @[system.scala 40:16]
  wire  rules_3_io_nT_out_1; // @[system.scala 40:16]
  wire  rules_3_io_nT_out_2; // @[system.scala 40:16]
  wire  rules_3_io_nC_in_0; // @[system.scala 40:16]
  wire  rules_3_io_nC_in_1; // @[system.scala 40:16]
  wire  rules_3_io_nC_in_2; // @[system.scala 40:16]
  wire  rules_3_io_nC_out_0; // @[system.scala 40:16]
  wire  rules_3_io_nC_out_1; // @[system.scala 40:16]
  wire  rules_3_io_nC_out_2; // @[system.scala 40:16]
  wire  rules_3_io_nE_in_0; // @[system.scala 40:16]
  wire  rules_3_io_nE_in_1; // @[system.scala 40:16]
  wire  rules_3_io_nE_in_2; // @[system.scala 40:16]
  wire  rules_3_io_nE_out_0; // @[system.scala 40:16]
  wire  rules_3_io_nE_out_1; // @[system.scala 40:16]
  wire  rules_3_io_nE_out_2; // @[system.scala 40:16]
  wire  rules_4_io_en_r; // @[system.scala 43:16]
  wire  rules_4_io_x_in; // @[system.scala 43:16]
  wire  rules_4_io_x_out; // @[system.scala 43:16]
  wire  rules_4_io_nI_in_0; // @[system.scala 43:16]
  wire  rules_4_io_nI_in_1; // @[system.scala 43:16]
  wire  rules_4_io_nI_in_2; // @[system.scala 43:16]
  wire  rules_4_io_nI_out_0; // @[system.scala 43:16]
  wire  rules_4_io_nI_out_1; // @[system.scala 43:16]
  wire  rules_4_io_nI_out_2; // @[system.scala 43:16]
  wire  rules_4_io_nT_in_0; // @[system.scala 43:16]
  wire  rules_4_io_nT_in_1; // @[system.scala 43:16]
  wire  rules_4_io_nT_in_2; // @[system.scala 43:16]
  wire  rules_4_io_nT_out_0; // @[system.scala 43:16]
  wire  rules_4_io_nT_out_1; // @[system.scala 43:16]
  wire  rules_4_io_nT_out_2; // @[system.scala 43:16]
  wire  rules_4_io_nC_in_0; // @[system.scala 43:16]
  wire  rules_4_io_nC_in_1; // @[system.scala 43:16]
  wire  rules_4_io_nC_in_2; // @[system.scala 43:16]
  wire  rules_4_io_nC_out_0; // @[system.scala 43:16]
  wire  rules_4_io_nC_out_1; // @[system.scala 43:16]
  wire  rules_4_io_nC_out_2; // @[system.scala 43:16]
  wire  rules_4_io_nE_in_0; // @[system.scala 43:16]
  wire  rules_4_io_nE_in_1; // @[system.scala 43:16]
  wire  rules_4_io_nE_in_2; // @[system.scala 43:16]
  wire  rules_4_io_nE_out_0; // @[system.scala 43:16]
  wire  rules_4_io_nE_out_1; // @[system.scala 43:16]
  wire  rules_4_io_nE_out_2; // @[system.scala 43:16]
  wire  rules_5_io_en_r; // @[system.scala 43:16]
  wire  rules_5_io_x_in; // @[system.scala 43:16]
  wire  rules_5_io_x_out; // @[system.scala 43:16]
  wire  rules_5_io_nI_in_0; // @[system.scala 43:16]
  wire  rules_5_io_nI_in_1; // @[system.scala 43:16]
  wire  rules_5_io_nI_in_2; // @[system.scala 43:16]
  wire  rules_5_io_nI_out_0; // @[system.scala 43:16]
  wire  rules_5_io_nI_out_1; // @[system.scala 43:16]
  wire  rules_5_io_nI_out_2; // @[system.scala 43:16]
  wire  rules_5_io_nT_in_0; // @[system.scala 43:16]
  wire  rules_5_io_nT_in_1; // @[system.scala 43:16]
  wire  rules_5_io_nT_in_2; // @[system.scala 43:16]
  wire  rules_5_io_nT_out_0; // @[system.scala 43:16]
  wire  rules_5_io_nT_out_1; // @[system.scala 43:16]
  wire  rules_5_io_nT_out_2; // @[system.scala 43:16]
  wire  rules_5_io_nC_in_0; // @[system.scala 43:16]
  wire  rules_5_io_nC_in_1; // @[system.scala 43:16]
  wire  rules_5_io_nC_in_2; // @[system.scala 43:16]
  wire  rules_5_io_nC_out_0; // @[system.scala 43:16]
  wire  rules_5_io_nC_out_1; // @[system.scala 43:16]
  wire  rules_5_io_nC_out_2; // @[system.scala 43:16]
  wire  rules_5_io_nE_in_0; // @[system.scala 43:16]
  wire  rules_5_io_nE_in_1; // @[system.scala 43:16]
  wire  rules_5_io_nE_in_2; // @[system.scala 43:16]
  wire  rules_5_io_nE_out_0; // @[system.scala 43:16]
  wire  rules_5_io_nE_out_1; // @[system.scala 43:16]
  wire  rules_5_io_nE_out_2; // @[system.scala 43:16]
  wire  rules_6_io_en_r; // @[system.scala 46:16]
  wire  rules_6_io_x_in; // @[system.scala 46:16]
  wire  rules_6_io_x_out; // @[system.scala 46:16]
  wire  rules_6_io_nI_in_0; // @[system.scala 46:16]
  wire  rules_6_io_nI_in_1; // @[system.scala 46:16]
  wire  rules_6_io_nI_in_2; // @[system.scala 46:16]
  wire  rules_6_io_nI_out_0; // @[system.scala 46:16]
  wire  rules_6_io_nI_out_1; // @[system.scala 46:16]
  wire  rules_6_io_nI_out_2; // @[system.scala 46:16]
  wire  rules_6_io_nT_in_0; // @[system.scala 46:16]
  wire  rules_6_io_nT_in_1; // @[system.scala 46:16]
  wire  rules_6_io_nT_in_2; // @[system.scala 46:16]
  wire  rules_6_io_nT_out_0; // @[system.scala 46:16]
  wire  rules_6_io_nT_out_1; // @[system.scala 46:16]
  wire  rules_6_io_nT_out_2; // @[system.scala 46:16]
  wire  rules_6_io_nC_in_0; // @[system.scala 46:16]
  wire  rules_6_io_nC_in_1; // @[system.scala 46:16]
  wire  rules_6_io_nC_in_2; // @[system.scala 46:16]
  wire  rules_6_io_nC_out_0; // @[system.scala 46:16]
  wire  rules_6_io_nC_out_1; // @[system.scala 46:16]
  wire  rules_6_io_nC_out_2; // @[system.scala 46:16]
  wire  rules_6_io_nE_in_0; // @[system.scala 46:16]
  wire  rules_6_io_nE_in_1; // @[system.scala 46:16]
  wire  rules_6_io_nE_in_2; // @[system.scala 46:16]
  wire  rules_6_io_nE_out_0; // @[system.scala 46:16]
  wire  rules_6_io_nE_out_1; // @[system.scala 46:16]
  wire  rules_6_io_nE_out_2; // @[system.scala 46:16]
  wire  rules_7_io_en_r; // @[system.scala 46:16]
  wire  rules_7_io_x_in; // @[system.scala 46:16]
  wire  rules_7_io_x_out; // @[system.scala 46:16]
  wire  rules_7_io_nI_in_0; // @[system.scala 46:16]
  wire  rules_7_io_nI_in_1; // @[system.scala 46:16]
  wire  rules_7_io_nI_in_2; // @[system.scala 46:16]
  wire  rules_7_io_nI_out_0; // @[system.scala 46:16]
  wire  rules_7_io_nI_out_1; // @[system.scala 46:16]
  wire  rules_7_io_nI_out_2; // @[system.scala 46:16]
  wire  rules_7_io_nT_in_0; // @[system.scala 46:16]
  wire  rules_7_io_nT_in_1; // @[system.scala 46:16]
  wire  rules_7_io_nT_in_2; // @[system.scala 46:16]
  wire  rules_7_io_nT_out_0; // @[system.scala 46:16]
  wire  rules_7_io_nT_out_1; // @[system.scala 46:16]
  wire  rules_7_io_nT_out_2; // @[system.scala 46:16]
  wire  rules_7_io_nC_in_0; // @[system.scala 46:16]
  wire  rules_7_io_nC_in_1; // @[system.scala 46:16]
  wire  rules_7_io_nC_in_2; // @[system.scala 46:16]
  wire  rules_7_io_nC_out_0; // @[system.scala 46:16]
  wire  rules_7_io_nC_out_1; // @[system.scala 46:16]
  wire  rules_7_io_nC_out_2; // @[system.scala 46:16]
  wire  rules_7_io_nE_in_0; // @[system.scala 46:16]
  wire  rules_7_io_nE_in_1; // @[system.scala 46:16]
  wire  rules_7_io_nE_in_2; // @[system.scala 46:16]
  wire  rules_7_io_nE_out_0; // @[system.scala 46:16]
  wire  rules_7_io_nE_out_1; // @[system.scala 46:16]
  wire  rules_7_io_nE_out_2; // @[system.scala 46:16]
  wire  rules_8_io_x_in; // @[system.scala 48:16]
  wire  rules_8_io_x_out; // @[system.scala 48:16]
  wire  rules_8_io_nI_in_0; // @[system.scala 48:16]
  wire  rules_8_io_nI_in_1; // @[system.scala 48:16]
  wire  rules_8_io_nI_in_2; // @[system.scala 48:16]
  wire  rules_8_io_nI_out_0; // @[system.scala 48:16]
  wire  rules_8_io_nI_out_1; // @[system.scala 48:16]
  wire  rules_8_io_nI_out_2; // @[system.scala 48:16]
  wire  rules_8_io_nT_in_0; // @[system.scala 48:16]
  wire  rules_8_io_nT_in_1; // @[system.scala 48:16]
  wire  rules_8_io_nT_in_2; // @[system.scala 48:16]
  wire  rules_8_io_nT_out_0; // @[system.scala 48:16]
  wire  rules_8_io_nT_out_1; // @[system.scala 48:16]
  wire  rules_8_io_nT_out_2; // @[system.scala 48:16]
  wire  rules_8_io_nC_in_0; // @[system.scala 48:16]
  wire  rules_8_io_nC_in_1; // @[system.scala 48:16]
  wire  rules_8_io_nC_in_2; // @[system.scala 48:16]
  wire  rules_8_io_nC_out_0; // @[system.scala 48:16]
  wire  rules_8_io_nC_out_1; // @[system.scala 48:16]
  wire  rules_8_io_nC_out_2; // @[system.scala 48:16]
  wire  rules_8_io_nE_in_0; // @[system.scala 48:16]
  wire  rules_8_io_nE_in_1; // @[system.scala 48:16]
  wire  rules_8_io_nE_in_2; // @[system.scala 48:16]
  wire  rules_8_io_nE_out_0; // @[system.scala 48:16]
  wire  rules_8_io_nE_out_1; // @[system.scala 48:16]
  wire  rules_8_io_nE_out_2; // @[system.scala 48:16]
  wire  rules_9_io_en_r; // @[system.scala 49:16]
  wire  rules_9_io_x_in; // @[system.scala 49:16]
  wire  rules_9_io_x_out; // @[system.scala 49:16]
  wire  rules_9_io_nI_in_0; // @[system.scala 49:16]
  wire  rules_9_io_nI_in_1; // @[system.scala 49:16]
  wire  rules_9_io_nI_in_2; // @[system.scala 49:16]
  wire  rules_9_io_nI_out_0; // @[system.scala 49:16]
  wire  rules_9_io_nI_out_1; // @[system.scala 49:16]
  wire  rules_9_io_nI_out_2; // @[system.scala 49:16]
  wire  rules_9_io_nT_in_0; // @[system.scala 49:16]
  wire  rules_9_io_nT_in_1; // @[system.scala 49:16]
  wire  rules_9_io_nT_in_2; // @[system.scala 49:16]
  wire  rules_9_io_nT_out_0; // @[system.scala 49:16]
  wire  rules_9_io_nT_out_1; // @[system.scala 49:16]
  wire  rules_9_io_nT_out_2; // @[system.scala 49:16]
  wire  rules_9_io_nC_in_0; // @[system.scala 49:16]
  wire  rules_9_io_nC_in_1; // @[system.scala 49:16]
  wire  rules_9_io_nC_in_2; // @[system.scala 49:16]
  wire  rules_9_io_nC_out_0; // @[system.scala 49:16]
  wire  rules_9_io_nC_out_1; // @[system.scala 49:16]
  wire  rules_9_io_nC_out_2; // @[system.scala 49:16]
  wire  rules_9_io_nE_in_0; // @[system.scala 49:16]
  wire  rules_9_io_nE_in_1; // @[system.scala 49:16]
  wire  rules_9_io_nE_in_2; // @[system.scala 49:16]
  wire  rules_9_io_nE_out_0; // @[system.scala 49:16]
  wire  rules_9_io_nE_out_1; // @[system.scala 49:16]
  wire  rules_9_io_nE_out_2; // @[system.scala 49:16]
  reg  x_reg; // @[system.scala 15:20]
  reg  nI_reg_0; // @[system.scala 18:21]
  reg  nI_reg_1; // @[system.scala 18:21]
  reg  nI_reg_2; // @[system.scala 18:21]
  reg  nT_reg_0; // @[system.scala 21:21]
  reg  nT_reg_1; // @[system.scala 21:21]
  reg  nT_reg_2; // @[system.scala 21:21]
  reg  nC_reg_0; // @[system.scala 24:21]
  reg  nC_reg_1; // @[system.scala 24:21]
  reg  nC_reg_2; // @[system.scala 24:21]
  reg  nE_reg_0; // @[system.scala 27:21]
  reg  nE_reg_1; // @[system.scala 27:21]
  reg  nE_reg_2; // @[system.scala 27:21]
  wire  _T = io_en_a == 4'h0; // @[system.scala 56:27]
  wire  _GEN_0 = _T ? rules_0_io_x_out : x_reg; // @[system.scala 15:20 57:21 58:7]
  wire  _GEN_1 = _T ? rules_0_io_nI_out_0 : nI_reg_0; // @[system.scala 18:21 57:21 59:8]
  wire  _GEN_2 = _T ? rules_0_io_nI_out_1 : nI_reg_1; // @[system.scala 18:21 57:21 59:8]
  wire  _GEN_3 = _T ? rules_0_io_nI_out_2 : nI_reg_2; // @[system.scala 18:21 57:21 59:8]
  wire  _GEN_4 = _T ? rules_0_io_nT_out_0 : nT_reg_0; // @[system.scala 21:21 57:21 60:8]
  wire  _GEN_5 = _T ? rules_0_io_nT_out_1 : nT_reg_1; // @[system.scala 21:21 57:21 60:8]
  wire  _GEN_6 = _T ? rules_0_io_nT_out_2 : nT_reg_2; // @[system.scala 21:21 57:21 60:8]
  wire  _GEN_7 = _T ? rules_0_io_nC_out_0 : nC_reg_0; // @[system.scala 24:21 57:21 61:8]
  wire  _GEN_8 = _T ? rules_0_io_nC_out_1 : nC_reg_1; // @[system.scala 24:21 57:21 61:8]
  wire  _GEN_9 = _T ? rules_0_io_nC_out_2 : nC_reg_2; // @[system.scala 24:21 57:21 61:8]
  wire  _GEN_10 = _T ? rules_0_io_nE_out_0 : nE_reg_0; // @[system.scala 27:21 57:21 62:8]
  wire  _GEN_11 = _T ? rules_0_io_nE_out_1 : nE_reg_1; // @[system.scala 27:21 57:21 62:8]
  wire  _GEN_12 = _T ? rules_0_io_nE_out_2 : nE_reg_2; // @[system.scala 27:21 57:21 62:8]
  wire  _T_2 = io_en_a == 4'h1; // @[system.scala 56:27]
  wire  _GEN_13 = _T_2 ? rules_1_io_x_out : _GEN_0; // @[system.scala 57:21 58:7]
  wire  _GEN_14 = _T_2 ? rules_1_io_nI_out_0 : _GEN_1; // @[system.scala 57:21 59:8]
  wire  _GEN_15 = _T_2 ? rules_1_io_nI_out_1 : _GEN_2; // @[system.scala 57:21 59:8]
  wire  _GEN_16 = _T_2 ? rules_1_io_nI_out_2 : _GEN_3; // @[system.scala 57:21 59:8]
  wire  _GEN_17 = _T_2 ? rules_1_io_nT_out_0 : _GEN_4; // @[system.scala 57:21 60:8]
  wire  _GEN_18 = _T_2 ? rules_1_io_nT_out_1 : _GEN_5; // @[system.scala 57:21 60:8]
  wire  _GEN_19 = _T_2 ? rules_1_io_nT_out_2 : _GEN_6; // @[system.scala 57:21 60:8]
  wire  _GEN_20 = _T_2 ? rules_1_io_nC_out_0 : _GEN_7; // @[system.scala 57:21 61:8]
  wire  _GEN_21 = _T_2 ? rules_1_io_nC_out_1 : _GEN_8; // @[system.scala 57:21 61:8]
  wire  _GEN_22 = _T_2 ? rules_1_io_nC_out_2 : _GEN_9; // @[system.scala 57:21 61:8]
  wire  _GEN_23 = _T_2 ? rules_1_io_nE_out_0 : _GEN_10; // @[system.scala 57:21 62:8]
  wire  _GEN_24 = _T_2 ? rules_1_io_nE_out_1 : _GEN_11; // @[system.scala 57:21 62:8]
  wire  _GEN_25 = _T_2 ? rules_1_io_nE_out_2 : _GEN_12; // @[system.scala 57:21 62:8]
  wire  _T_4 = io_en_a == 4'h2; // @[system.scala 56:27]
  wire  _GEN_26 = _T_4 ? rules_2_io_x_out : _GEN_13; // @[system.scala 57:21 58:7]
  wire  _GEN_27 = _T_4 ? rules_2_io_nI_out_0 : _GEN_14; // @[system.scala 57:21 59:8]
  wire  _GEN_28 = _T_4 ? rules_2_io_nI_out_1 : _GEN_15; // @[system.scala 57:21 59:8]
  wire  _GEN_29 = _T_4 ? rules_2_io_nI_out_2 : _GEN_16; // @[system.scala 57:21 59:8]
  wire  _GEN_30 = _T_4 ? rules_2_io_nT_out_0 : _GEN_17; // @[system.scala 57:21 60:8]
  wire  _GEN_31 = _T_4 ? rules_2_io_nT_out_1 : _GEN_18; // @[system.scala 57:21 60:8]
  wire  _GEN_32 = _T_4 ? rules_2_io_nT_out_2 : _GEN_19; // @[system.scala 57:21 60:8]
  wire  _GEN_33 = _T_4 ? rules_2_io_nC_out_0 : _GEN_20; // @[system.scala 57:21 61:8]
  wire  _GEN_34 = _T_4 ? rules_2_io_nC_out_1 : _GEN_21; // @[system.scala 57:21 61:8]
  wire  _GEN_35 = _T_4 ? rules_2_io_nC_out_2 : _GEN_22; // @[system.scala 57:21 61:8]
  wire  _GEN_36 = _T_4 ? rules_2_io_nE_out_0 : _GEN_23; // @[system.scala 57:21 62:8]
  wire  _GEN_37 = _T_4 ? rules_2_io_nE_out_1 : _GEN_24; // @[system.scala 57:21 62:8]
  wire  _GEN_38 = _T_4 ? rules_2_io_nE_out_2 : _GEN_25; // @[system.scala 57:21 62:8]
  wire  _T_6 = io_en_a == 4'h3; // @[system.scala 56:27]
  wire  _GEN_39 = _T_6 ? rules_3_io_x_out : _GEN_26; // @[system.scala 57:21 58:7]
  wire  _GEN_40 = _T_6 ? rules_3_io_nI_out_0 : _GEN_27; // @[system.scala 57:21 59:8]
  wire  _GEN_41 = _T_6 ? rules_3_io_nI_out_1 : _GEN_28; // @[system.scala 57:21 59:8]
  wire  _GEN_42 = _T_6 ? rules_3_io_nI_out_2 : _GEN_29; // @[system.scala 57:21 59:8]
  wire  _GEN_43 = _T_6 ? rules_3_io_nT_out_0 : _GEN_30; // @[system.scala 57:21 60:8]
  wire  _GEN_44 = _T_6 ? rules_3_io_nT_out_1 : _GEN_31; // @[system.scala 57:21 60:8]
  wire  _GEN_45 = _T_6 ? rules_3_io_nT_out_2 : _GEN_32; // @[system.scala 57:21 60:8]
  wire  _GEN_46 = _T_6 ? rules_3_io_nC_out_0 : _GEN_33; // @[system.scala 57:21 61:8]
  wire  _GEN_47 = _T_6 ? rules_3_io_nC_out_1 : _GEN_34; // @[system.scala 57:21 61:8]
  wire  _GEN_48 = _T_6 ? rules_3_io_nC_out_2 : _GEN_35; // @[system.scala 57:21 61:8]
  wire  _GEN_49 = _T_6 ? rules_3_io_nE_out_0 : _GEN_36; // @[system.scala 57:21 62:8]
  wire  _GEN_50 = _T_6 ? rules_3_io_nE_out_1 : _GEN_37; // @[system.scala 57:21 62:8]
  wire  _GEN_51 = _T_6 ? rules_3_io_nE_out_2 : _GEN_38; // @[system.scala 57:21 62:8]
  wire  _T_8 = io_en_a == 4'h4; // @[system.scala 56:27]
  wire  _GEN_52 = _T_8 ? rules_4_io_x_out : _GEN_39; // @[system.scala 57:21 58:7]
  wire  _GEN_53 = _T_8 ? rules_4_io_nI_out_0 : _GEN_40; // @[system.scala 57:21 59:8]
  wire  _GEN_54 = _T_8 ? rules_4_io_nI_out_1 : _GEN_41; // @[system.scala 57:21 59:8]
  wire  _GEN_55 = _T_8 ? rules_4_io_nI_out_2 : _GEN_42; // @[system.scala 57:21 59:8]
  wire  _GEN_56 = _T_8 ? rules_4_io_nT_out_0 : _GEN_43; // @[system.scala 57:21 60:8]
  wire  _GEN_57 = _T_8 ? rules_4_io_nT_out_1 : _GEN_44; // @[system.scala 57:21 60:8]
  wire  _GEN_58 = _T_8 ? rules_4_io_nT_out_2 : _GEN_45; // @[system.scala 57:21 60:8]
  wire  _GEN_59 = _T_8 ? rules_4_io_nC_out_0 : _GEN_46; // @[system.scala 57:21 61:8]
  wire  _GEN_60 = _T_8 ? rules_4_io_nC_out_1 : _GEN_47; // @[system.scala 57:21 61:8]
  wire  _GEN_61 = _T_8 ? rules_4_io_nC_out_2 : _GEN_48; // @[system.scala 57:21 61:8]
  wire  _GEN_62 = _T_8 ? rules_4_io_nE_out_0 : _GEN_49; // @[system.scala 57:21 62:8]
  wire  _GEN_63 = _T_8 ? rules_4_io_nE_out_1 : _GEN_50; // @[system.scala 57:21 62:8]
  wire  _GEN_64 = _T_8 ? rules_4_io_nE_out_2 : _GEN_51; // @[system.scala 57:21 62:8]
  wire  _T_10 = io_en_a == 4'h5; // @[system.scala 56:27]
  wire  _GEN_65 = _T_10 ? rules_5_io_x_out : _GEN_52; // @[system.scala 57:21 58:7]
  wire  _GEN_66 = _T_10 ? rules_5_io_nI_out_0 : _GEN_53; // @[system.scala 57:21 59:8]
  wire  _GEN_67 = _T_10 ? rules_5_io_nI_out_1 : _GEN_54; // @[system.scala 57:21 59:8]
  wire  _GEN_68 = _T_10 ? rules_5_io_nI_out_2 : _GEN_55; // @[system.scala 57:21 59:8]
  wire  _GEN_69 = _T_10 ? rules_5_io_nT_out_0 : _GEN_56; // @[system.scala 57:21 60:8]
  wire  _GEN_70 = _T_10 ? rules_5_io_nT_out_1 : _GEN_57; // @[system.scala 57:21 60:8]
  wire  _GEN_71 = _T_10 ? rules_5_io_nT_out_2 : _GEN_58; // @[system.scala 57:21 60:8]
  wire  _GEN_72 = _T_10 ? rules_5_io_nC_out_0 : _GEN_59; // @[system.scala 57:21 61:8]
  wire  _GEN_73 = _T_10 ? rules_5_io_nC_out_1 : _GEN_60; // @[system.scala 57:21 61:8]
  wire  _GEN_74 = _T_10 ? rules_5_io_nC_out_2 : _GEN_61; // @[system.scala 57:21 61:8]
  wire  _GEN_75 = _T_10 ? rules_5_io_nE_out_0 : _GEN_62; // @[system.scala 57:21 62:8]
  wire  _GEN_76 = _T_10 ? rules_5_io_nE_out_1 : _GEN_63; // @[system.scala 57:21 62:8]
  wire  _GEN_77 = _T_10 ? rules_5_io_nE_out_2 : _GEN_64; // @[system.scala 57:21 62:8]
  wire  _T_12 = io_en_a == 4'h6; // @[system.scala 56:27]
  wire  _GEN_78 = _T_12 ? rules_6_io_x_out : _GEN_65; // @[system.scala 57:21 58:7]
  wire  _GEN_79 = _T_12 ? rules_6_io_nI_out_0 : _GEN_66; // @[system.scala 57:21 59:8]
  wire  _GEN_80 = _T_12 ? rules_6_io_nI_out_1 : _GEN_67; // @[system.scala 57:21 59:8]
  wire  _GEN_81 = _T_12 ? rules_6_io_nI_out_2 : _GEN_68; // @[system.scala 57:21 59:8]
  wire  _GEN_82 = _T_12 ? rules_6_io_nT_out_0 : _GEN_69; // @[system.scala 57:21 60:8]
  wire  _GEN_83 = _T_12 ? rules_6_io_nT_out_1 : _GEN_70; // @[system.scala 57:21 60:8]
  wire  _GEN_84 = _T_12 ? rules_6_io_nT_out_2 : _GEN_71; // @[system.scala 57:21 60:8]
  wire  _GEN_85 = _T_12 ? rules_6_io_nC_out_0 : _GEN_72; // @[system.scala 57:21 61:8]
  wire  _GEN_86 = _T_12 ? rules_6_io_nC_out_1 : _GEN_73; // @[system.scala 57:21 61:8]
  wire  _GEN_87 = _T_12 ? rules_6_io_nC_out_2 : _GEN_74; // @[system.scala 57:21 61:8]
  wire  _GEN_88 = _T_12 ? rules_6_io_nE_out_0 : _GEN_75; // @[system.scala 57:21 62:8]
  wire  _GEN_89 = _T_12 ? rules_6_io_nE_out_1 : _GEN_76; // @[system.scala 57:21 62:8]
  wire  _GEN_90 = _T_12 ? rules_6_io_nE_out_2 : _GEN_77; // @[system.scala 57:21 62:8]
  wire  _T_14 = io_en_a == 4'h7; // @[system.scala 56:27]
  wire  _GEN_91 = _T_14 ? rules_7_io_x_out : _GEN_78; // @[system.scala 57:21 58:7]
  wire  _GEN_92 = _T_14 ? rules_7_io_nI_out_0 : _GEN_79; // @[system.scala 57:21 59:8]
  wire  _GEN_93 = _T_14 ? rules_7_io_nI_out_1 : _GEN_80; // @[system.scala 57:21 59:8]
  wire  _GEN_94 = _T_14 ? rules_7_io_nI_out_2 : _GEN_81; // @[system.scala 57:21 59:8]
  wire  _T_16 = io_en_a == 4'h8; // @[system.scala 56:27]
  wire  _GEN_104 = _T_16 ? rules_8_io_x_out : _GEN_91; // @[system.scala 57:21 58:7]
  wire  _GEN_105 = _T_16 ? rules_8_io_nI_out_0 : _GEN_92; // @[system.scala 57:21 59:8]
  wire  _GEN_106 = _T_16 ? rules_8_io_nI_out_1 : _GEN_93; // @[system.scala 57:21 59:8]
  wire  _GEN_107 = _T_16 ? rules_8_io_nI_out_2 : _GEN_94; // @[system.scala 57:21 59:8]
  wire  _T_18 = io_en_a == 4'h9; // @[system.scala 56:27]
  wire  _GEN_117 = _T_18 ? rules_9_io_x_out : _GEN_104; // @[system.scala 57:21 58:7]
  wire  _GEN_118 = _T_18 ? rules_9_io_nI_out_0 : _GEN_105; // @[system.scala 57:21 59:8]
  wire  _GEN_119 = _T_18 ? rules_9_io_nI_out_1 : _GEN_106; // @[system.scala 57:21 59:8]
  wire  _GEN_120 = _T_18 ? rules_9_io_nI_out_2 : _GEN_107; // @[system.scala 57:21 59:8]
  wire  _T_22 = ~nC_reg_1; // @[system.scala 75:24]
  wire  _T_27 = ~reset; // @[system.scala 75:7]
  wire  _T_32 = ~nC_reg_2; // @[system.scala 75:37]
  wire  _T_58 = ~nE_reg_1; // @[system.scala 80:24]
  wire  _T_68 = ~nE_reg_2; // @[system.scala 80:37]
  Try rules_0 ( // @[system.scala 37:16]
    .io_en_r(rules_0_io_en_r),
    .io_x_in(rules_0_io_x_in),
    .io_x_out(rules_0_io_x_out),
    .io_nI_in_0(rules_0_io_nI_in_0),
    .io_nI_in_1(rules_0_io_nI_in_1),
    .io_nI_in_2(rules_0_io_nI_in_2),
    .io_nI_out_0(rules_0_io_nI_out_0),
    .io_nI_out_1(rules_0_io_nI_out_1),
    .io_nI_out_2(rules_0_io_nI_out_2),
    .io_nT_in_0(rules_0_io_nT_in_0),
    .io_nT_in_1(rules_0_io_nT_in_1),
    .io_nT_in_2(rules_0_io_nT_in_2),
    .io_nT_out_0(rules_0_io_nT_out_0),
    .io_nT_out_1(rules_0_io_nT_out_1),
    .io_nT_out_2(rules_0_io_nT_out_2),
    .io_nC_in_0(rules_0_io_nC_in_0),
    .io_nC_in_1(rules_0_io_nC_in_1),
    .io_nC_in_2(rules_0_io_nC_in_2),
    .io_nC_out_0(rules_0_io_nC_out_0),
    .io_nC_out_1(rules_0_io_nC_out_1),
    .io_nC_out_2(rules_0_io_nC_out_2),
    .io_nE_in_0(rules_0_io_nE_in_0),
    .io_nE_in_1(rules_0_io_nE_in_1),
    .io_nE_in_2(rules_0_io_nE_in_2),
    .io_nE_out_0(rules_0_io_nE_out_0),
    .io_nE_out_1(rules_0_io_nE_out_1),
    .io_nE_out_2(rules_0_io_nE_out_2)
  );
  Try_1 rules_1 ( // @[system.scala 37:16]
    .io_en_r(rules_1_io_en_r),
    .io_x_in(rules_1_io_x_in),
    .io_x_out(rules_1_io_x_out),
    .io_nI_in_0(rules_1_io_nI_in_0),
    .io_nI_in_1(rules_1_io_nI_in_1),
    .io_nI_in_2(rules_1_io_nI_in_2),
    .io_nI_out_0(rules_1_io_nI_out_0),
    .io_nI_out_1(rules_1_io_nI_out_1),
    .io_nI_out_2(rules_1_io_nI_out_2),
    .io_nT_in_0(rules_1_io_nT_in_0),
    .io_nT_in_1(rules_1_io_nT_in_1),
    .io_nT_in_2(rules_1_io_nT_in_2),
    .io_nT_out_0(rules_1_io_nT_out_0),
    .io_nT_out_1(rules_1_io_nT_out_1),
    .io_nT_out_2(rules_1_io_nT_out_2),
    .io_nC_in_0(rules_1_io_nC_in_0),
    .io_nC_in_1(rules_1_io_nC_in_1),
    .io_nC_in_2(rules_1_io_nC_in_2),
    .io_nC_out_0(rules_1_io_nC_out_0),
    .io_nC_out_1(rules_1_io_nC_out_1),
    .io_nC_out_2(rules_1_io_nC_out_2),
    .io_nE_in_0(rules_1_io_nE_in_0),
    .io_nE_in_1(rules_1_io_nE_in_1),
    .io_nE_in_2(rules_1_io_nE_in_2),
    .io_nE_out_0(rules_1_io_nE_out_0),
    .io_nE_out_1(rules_1_io_nE_out_1),
    .io_nE_out_2(rules_1_io_nE_out_2)
  );
  Crit rules_2 ( // @[system.scala 40:16]
    .io_en_r(rules_2_io_en_r),
    .io_x_in(rules_2_io_x_in),
    .io_x_out(rules_2_io_x_out),
    .io_nI_in_0(rules_2_io_nI_in_0),
    .io_nI_in_1(rules_2_io_nI_in_1),
    .io_nI_in_2(rules_2_io_nI_in_2),
    .io_nI_out_0(rules_2_io_nI_out_0),
    .io_nI_out_1(rules_2_io_nI_out_1),
    .io_nI_out_2(rules_2_io_nI_out_2),
    .io_nT_in_0(rules_2_io_nT_in_0),
    .io_nT_in_1(rules_2_io_nT_in_1),
    .io_nT_in_2(rules_2_io_nT_in_2),
    .io_nT_out_0(rules_2_io_nT_out_0),
    .io_nT_out_1(rules_2_io_nT_out_1),
    .io_nT_out_2(rules_2_io_nT_out_2),
    .io_nC_in_0(rules_2_io_nC_in_0),
    .io_nC_in_1(rules_2_io_nC_in_1),
    .io_nC_in_2(rules_2_io_nC_in_2),
    .io_nC_out_0(rules_2_io_nC_out_0),
    .io_nC_out_1(rules_2_io_nC_out_1),
    .io_nC_out_2(rules_2_io_nC_out_2),
    .io_nE_in_0(rules_2_io_nE_in_0),
    .io_nE_in_1(rules_2_io_nE_in_1),
    .io_nE_in_2(rules_2_io_nE_in_2),
    .io_nE_out_0(rules_2_io_nE_out_0),
    .io_nE_out_1(rules_2_io_nE_out_1),
    .io_nE_out_2(rules_2_io_nE_out_2)
  );
  Crit_1 rules_3 ( // @[system.scala 40:16]
    .io_en_r(rules_3_io_en_r),
    .io_x_in(rules_3_io_x_in),
    .io_x_out(rules_3_io_x_out),
    .io_nI_in_0(rules_3_io_nI_in_0),
    .io_nI_in_1(rules_3_io_nI_in_1),
    .io_nI_in_2(rules_3_io_nI_in_2),
    .io_nI_out_0(rules_3_io_nI_out_0),
    .io_nI_out_1(rules_3_io_nI_out_1),
    .io_nI_out_2(rules_3_io_nI_out_2),
    .io_nT_in_0(rules_3_io_nT_in_0),
    .io_nT_in_1(rules_3_io_nT_in_1),
    .io_nT_in_2(rules_3_io_nT_in_2),
    .io_nT_out_0(rules_3_io_nT_out_0),
    .io_nT_out_1(rules_3_io_nT_out_1),
    .io_nT_out_2(rules_3_io_nT_out_2),
    .io_nC_in_0(rules_3_io_nC_in_0),
    .io_nC_in_1(rules_3_io_nC_in_1),
    .io_nC_in_2(rules_3_io_nC_in_2),
    .io_nC_out_0(rules_3_io_nC_out_0),
    .io_nC_out_1(rules_3_io_nC_out_1),
    .io_nC_out_2(rules_3_io_nC_out_2),
    .io_nE_in_0(rules_3_io_nE_in_0),
    .io_nE_in_1(rules_3_io_nE_in_1),
    .io_nE_in_2(rules_3_io_nE_in_2),
    .io_nE_out_0(rules_3_io_nE_out_0),
    .io_nE_out_1(rules_3_io_nE_out_1),
    .io_nE_out_2(rules_3_io_nE_out_2)
  );
  Exit rules_4 ( // @[system.scala 43:16]
    .io_en_r(rules_4_io_en_r),
    .io_x_in(rules_4_io_x_in),
    .io_x_out(rules_4_io_x_out),
    .io_nI_in_0(rules_4_io_nI_in_0),
    .io_nI_in_1(rules_4_io_nI_in_1),
    .io_nI_in_2(rules_4_io_nI_in_2),
    .io_nI_out_0(rules_4_io_nI_out_0),
    .io_nI_out_1(rules_4_io_nI_out_1),
    .io_nI_out_2(rules_4_io_nI_out_2),
    .io_nT_in_0(rules_4_io_nT_in_0),
    .io_nT_in_1(rules_4_io_nT_in_1),
    .io_nT_in_2(rules_4_io_nT_in_2),
    .io_nT_out_0(rules_4_io_nT_out_0),
    .io_nT_out_1(rules_4_io_nT_out_1),
    .io_nT_out_2(rules_4_io_nT_out_2),
    .io_nC_in_0(rules_4_io_nC_in_0),
    .io_nC_in_1(rules_4_io_nC_in_1),
    .io_nC_in_2(rules_4_io_nC_in_2),
    .io_nC_out_0(rules_4_io_nC_out_0),
    .io_nC_out_1(rules_4_io_nC_out_1),
    .io_nC_out_2(rules_4_io_nC_out_2),
    .io_nE_in_0(rules_4_io_nE_in_0),
    .io_nE_in_1(rules_4_io_nE_in_1),
    .io_nE_in_2(rules_4_io_nE_in_2),
    .io_nE_out_0(rules_4_io_nE_out_0),
    .io_nE_out_1(rules_4_io_nE_out_1),
    .io_nE_out_2(rules_4_io_nE_out_2)
  );
  Exit_1 rules_5 ( // @[system.scala 43:16]
    .io_en_r(rules_5_io_en_r),
    .io_x_in(rules_5_io_x_in),
    .io_x_out(rules_5_io_x_out),
    .io_nI_in_0(rules_5_io_nI_in_0),
    .io_nI_in_1(rules_5_io_nI_in_1),
    .io_nI_in_2(rules_5_io_nI_in_2),
    .io_nI_out_0(rules_5_io_nI_out_0),
    .io_nI_out_1(rules_5_io_nI_out_1),
    .io_nI_out_2(rules_5_io_nI_out_2),
    .io_nT_in_0(rules_5_io_nT_in_0),
    .io_nT_in_1(rules_5_io_nT_in_1),
    .io_nT_in_2(rules_5_io_nT_in_2),
    .io_nT_out_0(rules_5_io_nT_out_0),
    .io_nT_out_1(rules_5_io_nT_out_1),
    .io_nT_out_2(rules_5_io_nT_out_2),
    .io_nC_in_0(rules_5_io_nC_in_0),
    .io_nC_in_1(rules_5_io_nC_in_1),
    .io_nC_in_2(rules_5_io_nC_in_2),
    .io_nC_out_0(rules_5_io_nC_out_0),
    .io_nC_out_1(rules_5_io_nC_out_1),
    .io_nC_out_2(rules_5_io_nC_out_2),
    .io_nE_in_0(rules_5_io_nE_in_0),
    .io_nE_in_1(rules_5_io_nE_in_1),
    .io_nE_in_2(rules_5_io_nE_in_2),
    .io_nE_out_0(rules_5_io_nE_out_0),
    .io_nE_out_1(rules_5_io_nE_out_1),
    .io_nE_out_2(rules_5_io_nE_out_2)
  );
  Idle rules_6 ( // @[system.scala 46:16]
    .io_en_r(rules_6_io_en_r),
    .io_x_in(rules_6_io_x_in),
    .io_x_out(rules_6_io_x_out),
    .io_nI_in_0(rules_6_io_nI_in_0),
    .io_nI_in_1(rules_6_io_nI_in_1),
    .io_nI_in_2(rules_6_io_nI_in_2),
    .io_nI_out_0(rules_6_io_nI_out_0),
    .io_nI_out_1(rules_6_io_nI_out_1),
    .io_nI_out_2(rules_6_io_nI_out_2),
    .io_nT_in_0(rules_6_io_nT_in_0),
    .io_nT_in_1(rules_6_io_nT_in_1),
    .io_nT_in_2(rules_6_io_nT_in_2),
    .io_nT_out_0(rules_6_io_nT_out_0),
    .io_nT_out_1(rules_6_io_nT_out_1),
    .io_nT_out_2(rules_6_io_nT_out_2),
    .io_nC_in_0(rules_6_io_nC_in_0),
    .io_nC_in_1(rules_6_io_nC_in_1),
    .io_nC_in_2(rules_6_io_nC_in_2),
    .io_nC_out_0(rules_6_io_nC_out_0),
    .io_nC_out_1(rules_6_io_nC_out_1),
    .io_nC_out_2(rules_6_io_nC_out_2),
    .io_nE_in_0(rules_6_io_nE_in_0),
    .io_nE_in_1(rules_6_io_nE_in_1),
    .io_nE_in_2(rules_6_io_nE_in_2),
    .io_nE_out_0(rules_6_io_nE_out_0),
    .io_nE_out_1(rules_6_io_nE_out_1),
    .io_nE_out_2(rules_6_io_nE_out_2)
  );
  Idle_1 rules_7 ( // @[system.scala 46:16]
    .io_en_r(rules_7_io_en_r),
    .io_x_in(rules_7_io_x_in),
    .io_x_out(rules_7_io_x_out),
    .io_nI_in_0(rules_7_io_nI_in_0),
    .io_nI_in_1(rules_7_io_nI_in_1),
    .io_nI_in_2(rules_7_io_nI_in_2),
    .io_nI_out_0(rules_7_io_nI_out_0),
    .io_nI_out_1(rules_7_io_nI_out_1),
    .io_nI_out_2(rules_7_io_nI_out_2),
    .io_nT_in_0(rules_7_io_nT_in_0),
    .io_nT_in_1(rules_7_io_nT_in_1),
    .io_nT_in_2(rules_7_io_nT_in_2),
    .io_nT_out_0(rules_7_io_nT_out_0),
    .io_nT_out_1(rules_7_io_nT_out_1),
    .io_nT_out_2(rules_7_io_nT_out_2),
    .io_nC_in_0(rules_7_io_nC_in_0),
    .io_nC_in_1(rules_7_io_nC_in_1),
    .io_nC_in_2(rules_7_io_nC_in_2),
    .io_nC_out_0(rules_7_io_nC_out_0),
    .io_nC_out_1(rules_7_io_nC_out_1),
    .io_nC_out_2(rules_7_io_nC_out_2),
    .io_nE_in_0(rules_7_io_nE_in_0),
    .io_nE_in_1(rules_7_io_nE_in_1),
    .io_nE_in_2(rules_7_io_nE_in_2),
    .io_nE_out_0(rules_7_io_nE_out_0),
    .io_nE_out_1(rules_7_io_nE_out_1),
    .io_nE_out_2(rules_7_io_nE_out_2)
  );
  Str_Idle rules_8 ( // @[system.scala 48:16]
    .io_x_in(rules_8_io_x_in),
    .io_x_out(rules_8_io_x_out),
    .io_nI_in_0(rules_8_io_nI_in_0),
    .io_nI_in_1(rules_8_io_nI_in_1),
    .io_nI_in_2(rules_8_io_nI_in_2),
    .io_nI_out_0(rules_8_io_nI_out_0),
    .io_nI_out_1(rules_8_io_nI_out_1),
    .io_nI_out_2(rules_8_io_nI_out_2),
    .io_nT_in_0(rules_8_io_nT_in_0),
    .io_nT_in_1(rules_8_io_nT_in_1),
    .io_nT_in_2(rules_8_io_nT_in_2),
    .io_nT_out_0(rules_8_io_nT_out_0),
    .io_nT_out_1(rules_8_io_nT_out_1),
    .io_nT_out_2(rules_8_io_nT_out_2),
    .io_nC_in_0(rules_8_io_nC_in_0),
    .io_nC_in_1(rules_8_io_nC_in_1),
    .io_nC_in_2(rules_8_io_nC_in_2),
    .io_nC_out_0(rules_8_io_nC_out_0),
    .io_nC_out_1(rules_8_io_nC_out_1),
    .io_nC_out_2(rules_8_io_nC_out_2),
    .io_nE_in_0(rules_8_io_nE_in_0),
    .io_nE_in_1(rules_8_io_nE_in_1),
    .io_nE_in_2(rules_8_io_nE_in_2),
    .io_nE_out_0(rules_8_io_nE_out_0),
    .io_nE_out_1(rules_8_io_nE_out_1),
    .io_nE_out_2(rules_8_io_nE_out_2)
  );
  Str_Crit rules_9 ( // @[system.scala 49:16]
    .io_en_r(rules_9_io_en_r),
    .io_x_in(rules_9_io_x_in),
    .io_x_out(rules_9_io_x_out),
    .io_nI_in_0(rules_9_io_nI_in_0),
    .io_nI_in_1(rules_9_io_nI_in_1),
    .io_nI_in_2(rules_9_io_nI_in_2),
    .io_nI_out_0(rules_9_io_nI_out_0),
    .io_nI_out_1(rules_9_io_nI_out_1),
    .io_nI_out_2(rules_9_io_nI_out_2),
    .io_nT_in_0(rules_9_io_nT_in_0),
    .io_nT_in_1(rules_9_io_nT_in_1),
    .io_nT_in_2(rules_9_io_nT_in_2),
    .io_nT_out_0(rules_9_io_nT_out_0),
    .io_nT_out_1(rules_9_io_nT_out_1),
    .io_nT_out_2(rules_9_io_nT_out_2),
    .io_nC_in_0(rules_9_io_nC_in_0),
    .io_nC_in_1(rules_9_io_nC_in_1),
    .io_nC_in_2(rules_9_io_nC_in_2),
    .io_nC_out_0(rules_9_io_nC_out_0),
    .io_nC_out_1(rules_9_io_nC_out_1),
    .io_nC_out_2(rules_9_io_nC_out_2),
    .io_nE_in_0(rules_9_io_nE_in_0),
    .io_nE_in_1(rules_9_io_nE_in_1),
    .io_nE_in_2(rules_9_io_nE_in_2),
    .io_nE_out_0(rules_9_io_nE_out_0),
    .io_nE_out_1(rules_9_io_nE_out_1),
    .io_nE_out_2(rules_9_io_nE_out_2)
  );
  assign io_x_out = x_reg; // @[system.scala 16:9]
  assign io_nI_out_0 = nI_reg_0; // @[system.scala 19:10]
  assign io_nI_out_1 = nI_reg_1; // @[system.scala 19:10]
  assign io_nI_out_2 = nI_reg_2; // @[system.scala 19:10]
  assign io_nT_out_0 = nT_reg_0; // @[system.scala 22:10]
  assign io_nT_out_1 = nT_reg_1; // @[system.scala 22:10]
  assign io_nT_out_2 = nT_reg_2; // @[system.scala 22:10]
  assign io_nC_out_0 = nC_reg_0; // @[system.scala 25:10]
  assign io_nC_out_1 = nC_reg_1; // @[system.scala 25:10]
  assign io_nC_out_2 = nC_reg_2; // @[system.scala 25:10]
  assign io_nE_out_0 = nE_reg_0; // @[system.scala 28:10]
  assign io_nE_out_1 = nE_reg_1; // @[system.scala 28:10]
  assign io_nE_out_2 = nE_reg_2; // @[system.scala 28:10]
  assign rules_0_io_en_r = io_en_a == 4'h0; // @[system.scala 56:27]
  assign rules_0_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_0_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_0_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_0_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_0_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_0_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_0_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_0_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_0_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_0_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_0_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_0_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_0_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_1_io_en_r = io_en_a == 4'h1; // @[system.scala 56:27]
  assign rules_1_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_1_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_1_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_1_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_1_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_1_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_1_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_1_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_1_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_1_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_1_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_1_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_1_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_2_io_en_r = io_en_a == 4'h2; // @[system.scala 56:27]
  assign rules_2_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_2_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_2_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_2_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_2_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_2_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_2_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_2_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_2_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_2_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_2_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_2_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_2_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_3_io_en_r = io_en_a == 4'h3; // @[system.scala 56:27]
  assign rules_3_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_3_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_3_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_3_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_3_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_3_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_3_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_3_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_3_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_3_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_3_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_3_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_3_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_4_io_en_r = io_en_a == 4'h4; // @[system.scala 56:27]
  assign rules_4_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_4_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_4_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_4_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_4_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_4_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_4_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_4_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_4_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_4_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_4_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_4_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_4_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_5_io_en_r = io_en_a == 4'h5; // @[system.scala 56:27]
  assign rules_5_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_5_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_5_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_5_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_5_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_5_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_5_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_5_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_5_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_5_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_5_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_5_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_5_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_6_io_en_r = io_en_a == 4'h6; // @[system.scala 56:27]
  assign rules_6_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_6_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_6_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_6_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_6_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_6_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_6_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_6_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_6_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_6_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_6_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_6_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_6_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_7_io_en_r = io_en_a == 4'h7; // @[system.scala 56:27]
  assign rules_7_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_7_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_7_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_7_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_7_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_7_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_7_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_7_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_7_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_7_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_7_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_7_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_7_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_8_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_8_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_8_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_8_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_8_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_8_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_8_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_8_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_8_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_8_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_8_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_8_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_8_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  assign rules_9_io_en_r = io_en_a == 4'h9; // @[system.scala 56:27]
  assign rules_9_io_x_in = x_reg; // @[system.scala 51:18]
  assign rules_9_io_nI_in_0 = nI_reg_0; // @[system.scala 52:19]
  assign rules_9_io_nI_in_1 = nI_reg_1; // @[system.scala 52:19]
  assign rules_9_io_nI_in_2 = nI_reg_2; // @[system.scala 52:19]
  assign rules_9_io_nT_in_0 = nT_reg_0; // @[system.scala 53:19]
  assign rules_9_io_nT_in_1 = nT_reg_1; // @[system.scala 53:19]
  assign rules_9_io_nT_in_2 = nT_reg_2; // @[system.scala 53:19]
  assign rules_9_io_nC_in_0 = nC_reg_0; // @[system.scala 54:19]
  assign rules_9_io_nC_in_1 = nC_reg_1; // @[system.scala 54:19]
  assign rules_9_io_nC_in_2 = nC_reg_2; // @[system.scala 54:19]
  assign rules_9_io_nE_in_0 = nE_reg_0; // @[system.scala 55:19]
  assign rules_9_io_nE_in_1 = nE_reg_1; // @[system.scala 55:19]
  assign rules_9_io_nE_in_2 = nE_reg_2; // @[system.scala 55:19]
  always @(posedge clock) begin
    x_reg <= reset | _GEN_117; // @[system.scala 15:{20,20}]
    nI_reg_0 <= reset | _GEN_118; // @[system.scala 18:{21,21}]
    nI_reg_1 <= reset | _GEN_119; // @[system.scala 18:{21,21}]
    nI_reg_2 <= reset | _GEN_120; // @[system.scala 18:{21,21}]
    if (reset) begin // @[system.scala 21:21]
      nT_reg_0 <= 1'h0; // @[system.scala 21:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nT_reg_0 <= rules_9_io_nT_out_0; // @[system.scala 60:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nT_reg_0 <= rules_8_io_nT_out_0; // @[system.scala 60:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nT_reg_0 <= rules_7_io_nT_out_0; // @[system.scala 60:8]
    end else begin
      nT_reg_0 <= _GEN_82;
    end
    if (reset) begin // @[system.scala 21:21]
      nT_reg_1 <= 1'h0; // @[system.scala 21:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nT_reg_1 <= rules_9_io_nT_out_1; // @[system.scala 60:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nT_reg_1 <= rules_8_io_nT_out_1; // @[system.scala 60:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nT_reg_1 <= rules_7_io_nT_out_1; // @[system.scala 60:8]
    end else begin
      nT_reg_1 <= _GEN_83;
    end
    if (reset) begin // @[system.scala 21:21]
      nT_reg_2 <= 1'h0; // @[system.scala 21:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nT_reg_2 <= rules_9_io_nT_out_2; // @[system.scala 60:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nT_reg_2 <= rules_8_io_nT_out_2; // @[system.scala 60:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nT_reg_2 <= rules_7_io_nT_out_2; // @[system.scala 60:8]
    end else begin
      nT_reg_2 <= _GEN_84;
    end
    if (reset) begin // @[system.scala 24:21]
      nC_reg_0 <= 1'h0; // @[system.scala 24:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nC_reg_0 <= rules_9_io_nC_out_0; // @[system.scala 61:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nC_reg_0 <= rules_8_io_nC_out_0; // @[system.scala 61:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nC_reg_0 <= rules_7_io_nC_out_0; // @[system.scala 61:8]
    end else begin
      nC_reg_0 <= _GEN_85;
    end
    if (reset) begin // @[system.scala 24:21]
      nC_reg_1 <= 1'h0; // @[system.scala 24:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nC_reg_1 <= rules_9_io_nC_out_1; // @[system.scala 61:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nC_reg_1 <= rules_8_io_nC_out_1; // @[system.scala 61:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nC_reg_1 <= rules_7_io_nC_out_1; // @[system.scala 61:8]
    end else begin
      nC_reg_1 <= _GEN_86;
    end
    if (reset) begin // @[system.scala 24:21]
      nC_reg_2 <= 1'h0; // @[system.scala 24:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nC_reg_2 <= rules_9_io_nC_out_2; // @[system.scala 61:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nC_reg_2 <= rules_8_io_nC_out_2; // @[system.scala 61:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nC_reg_2 <= rules_7_io_nC_out_2; // @[system.scala 61:8]
    end else begin
      nC_reg_2 <= _GEN_87;
    end
    if (reset) begin // @[system.scala 27:21]
      nE_reg_0 <= 1'h0; // @[system.scala 27:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nE_reg_0 <= rules_9_io_nE_out_0; // @[system.scala 62:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nE_reg_0 <= rules_8_io_nE_out_0; // @[system.scala 62:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nE_reg_0 <= rules_7_io_nE_out_0; // @[system.scala 62:8]
    end else begin
      nE_reg_0 <= _GEN_88;
    end
    if (reset) begin // @[system.scala 27:21]
      nE_reg_1 <= 1'h0; // @[system.scala 27:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nE_reg_1 <= rules_9_io_nE_out_1; // @[system.scala 62:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nE_reg_1 <= rules_8_io_nE_out_1; // @[system.scala 62:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nE_reg_1 <= rules_7_io_nE_out_1; // @[system.scala 62:8]
    end else begin
      nE_reg_1 <= _GEN_89;
    end
    if (reset) begin // @[system.scala 27:21]
      nE_reg_2 <= 1'h0; // @[system.scala 27:21]
    end else if (_T_18) begin // @[system.scala 57:21]
      nE_reg_2 <= rules_9_io_nE_out_2; // @[system.scala 62:8]
    end else if (_T_16) begin // @[system.scala 57:21]
      nE_reg_2 <= rules_8_io_nE_out_2; // @[system.scala 62:8]
    end else if (_T_14) begin // @[system.scala 57:21]
      nE_reg_2 <= rules_7_io_nE_out_2; // @[system.scala 62:8]
    end else begin
      nE_reg_2 <= _GEN_90;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif

                initial begin
                    assume(reset==1);
                end

                  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 75:7]
    end
    //
    if (~reset) begin
      assert(~nC_reg_1 | ~nC_reg_2); // @[system.scala 75:7]
    end
    //
    if (~reset) begin
      assert(~nC_reg_2 | ~nC_reg_1); // @[system.scala 75:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 75:7]
    end
    //
    if (_T_27) begin
      assert(1'h1); // @[system.scala 80:7]
    end
    //
    if (_T_27) begin
      assert(~nE_reg_1 | ~nE_reg_2); // @[system.scala 80:7]
    end
    //
    if (_T_27) begin
      assert(~nE_reg_2 | ~nE_reg_1); // @[system.scala 80:7]
    end
    //
    if (_T_27) begin
      assert(1'h1); // @[system.scala 80:7]
    end
    //
    if (_T_27) begin
      assert(1'h1); // @[system.scala 85:7]
    end
    //
    if (_T_27) begin
      assert(_T_58 | _T_32); // @[system.scala 85:7]
    end
    //
    if (_T_27) begin
      assert(_T_68 | _T_22); // @[system.scala 85:7]
    end
    //
    if (_T_27) begin
      assert(1'h1); // @[system.scala 85:7]
    end
  end
endmodule
