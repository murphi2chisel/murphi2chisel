module Init(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_en_r ? 2'h0 : io_n_in_1; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_2 = io_en_r ? 2'h0 : io_n_in_2; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_3 = io_en_r ? 2'h0 : io_n_in_3; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_4 = io_en_r ? 2'h0 : io_n_in_4; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_5 = io_en_r ? 2'h0 : io_n_in_5; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_6 = io_en_r ? 2'h0 : io_n_in_6; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_7 = io_en_r ? 2'h0 : io_n_in_7; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_8 = io_en_r ? 2'h0 : io_n_in_8; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_9 = io_en_r ? 2'h0 : io_n_in_9; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_10 = io_en_r ? 2'h0 : io_n_in_10; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_11 = io_en_r ? 2'h0 : io_n_in_11; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_12 = io_en_r ? 2'h0 : io_n_in_12; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_13 = io_en_r ? 2'h0 : io_n_in_13; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_14 = io_en_r ? 2'h0 : io_n_in_14; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_15 = io_en_r ? 2'h0 : io_n_in_15; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_n_out_16 = io_en_r ? 2'h0 : io_n_in_16; // @[router.scala 5:14 7:13 node.scala 30:9]
  assign io_x_out = io_en_r | io_x_in; // @[router.scala 10:10 5:14 node.scala 31:9]
endmodule
module Try(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_1 == 2'h0 ? 2'h1 : io_n_in_1; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_en_r ? _GEN_0 : io_n_in_1; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_1(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_2 == 2'h0 ? 2'h1 : io_n_in_2; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_en_r ? _GEN_0 : io_n_in_2; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_2(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_3 == 2'h0 ? 2'h1 : io_n_in_3; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_en_r ? _GEN_0 : io_n_in_3; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_3(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_4 == 2'h0 ? 2'h1 : io_n_in_4; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_en_r ? _GEN_0 : io_n_in_4; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_4(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_5 == 2'h0 ? 2'h1 : io_n_in_5; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_en_r ? _GEN_0 : io_n_in_5; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_5(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_6 == 2'h0 ? 2'h1 : io_n_in_6; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_en_r ? _GEN_0 : io_n_in_6; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_6(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_7 == 2'h0 ? 2'h1 : io_n_in_7; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_en_r ? _GEN_0 : io_n_in_7; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_7(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_8 == 2'h0 ? 2'h1 : io_n_in_8; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_en_r ? _GEN_0 : io_n_in_8; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_8(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_9 == 2'h0 ? 2'h1 : io_n_in_9; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_en_r ? _GEN_0 : io_n_in_9; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_9(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_10 == 2'h0 ? 2'h1 : io_n_in_10; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_en_r ? _GEN_0 : io_n_in_10; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_10(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_11 == 2'h0 ? 2'h1 : io_n_in_11; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_en_r ? _GEN_0 : io_n_in_11; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_11(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_12 == 2'h0 ? 2'h1 : io_n_in_12; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_en_r ? _GEN_0 : io_n_in_12; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_12(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_13 == 2'h0 ? 2'h1 : io_n_in_13; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_en_r ? _GEN_0 : io_n_in_13; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_13(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_14 == 2'h0 ? 2'h1 : io_n_in_14; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_en_r ? _GEN_0 : io_n_in_14; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_14(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_15 == 2'h0 ? 2'h1 : io_n_in_15; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_en_r ? _GEN_0 : io_n_in_15; // @[router.scala 14:14 node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Try_15(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_16 == 2'h0 ? 2'h1 : io_n_in_16; // @[router.scala 15:23 16:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_en_r ? _GEN_0 : io_n_in_16; // @[router.scala 14:14 node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Crit(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_1 == 2'h1 & io_x_in ? 2'h2 : io_n_in_1; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_1 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_en_r ? _GEN_0 : io_n_in_1; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_1(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_2 == 2'h1 & io_x_in ? 2'h2 : io_n_in_2; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_2 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_en_r ? _GEN_0 : io_n_in_2; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_2(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_3 == 2'h1 & io_x_in ? 2'h2 : io_n_in_3; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_3 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_en_r ? _GEN_0 : io_n_in_3; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_3(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_4 == 2'h1 & io_x_in ? 2'h2 : io_n_in_4; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_4 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_en_r ? _GEN_0 : io_n_in_4; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_4(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_5 == 2'h1 & io_x_in ? 2'h2 : io_n_in_5; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_5 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_en_r ? _GEN_0 : io_n_in_5; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_5(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_6 == 2'h1 & io_x_in ? 2'h2 : io_n_in_6; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_6 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_en_r ? _GEN_0 : io_n_in_6; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_6(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_7 == 2'h1 & io_x_in ? 2'h2 : io_n_in_7; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_7 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_en_r ? _GEN_0 : io_n_in_7; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_7(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_8 == 2'h1 & io_x_in ? 2'h2 : io_n_in_8; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_8 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_en_r ? _GEN_0 : io_n_in_8; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_8(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_9 == 2'h1 & io_x_in ? 2'h2 : io_n_in_9; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_9 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_en_r ? _GEN_0 : io_n_in_9; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_9(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_10 == 2'h1 & io_x_in ? 2'h2 : io_n_in_10; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_10 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_en_r ? _GEN_0 : io_n_in_10; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_10(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_11 == 2'h1 & io_x_in ? 2'h2 : io_n_in_11; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_11 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_en_r ? _GEN_0 : io_n_in_11; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_11(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_12 == 2'h1 & io_x_in ? 2'h2 : io_n_in_12; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_12 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_en_r ? _GEN_0 : io_n_in_12; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_12(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_13 == 2'h1 & io_x_in ? 2'h2 : io_n_in_13; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_13 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_en_r ? _GEN_0 : io_n_in_13; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_13(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_14 == 2'h1 & io_x_in ? 2'h2 : io_n_in_14; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_14 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_en_r ? _GEN_0 : io_n_in_14; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_14(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_15 == 2'h1 & io_x_in ? 2'h2 : io_n_in_15; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_15 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_en_r ? _GEN_0 : io_n_in_15; // @[router.scala 21:14 node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Crit_15(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_16 == 2'h1 & io_x_in ? 2'h2 : io_n_in_16; // @[router.scala 22:45 23:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_16 == 2'h1 & io_x_in ? 1'h0 : io_x_in; // @[router.scala 22:45 24:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_en_r ? _GEN_0 : io_n_in_16; // @[router.scala 21:14 node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 21:14 node.scala 31:9]
endmodule
module Exit(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_1 == 2'h2 ? 2'h3 : io_n_in_1; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_en_r ? _GEN_0 : io_n_in_1; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_1(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_2 == 2'h2 ? 2'h3 : io_n_in_2; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_en_r ? _GEN_0 : io_n_in_2; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_2(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_3 == 2'h2 ? 2'h3 : io_n_in_3; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_en_r ? _GEN_0 : io_n_in_3; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_3(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_4 == 2'h2 ? 2'h3 : io_n_in_4; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_en_r ? _GEN_0 : io_n_in_4; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_4(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_5 == 2'h2 ? 2'h3 : io_n_in_5; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_en_r ? _GEN_0 : io_n_in_5; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_5(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_6 == 2'h2 ? 2'h3 : io_n_in_6; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_en_r ? _GEN_0 : io_n_in_6; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_6(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_7 == 2'h2 ? 2'h3 : io_n_in_7; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_en_r ? _GEN_0 : io_n_in_7; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_7(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_8 == 2'h2 ? 2'h3 : io_n_in_8; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_en_r ? _GEN_0 : io_n_in_8; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_8(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_9 == 2'h2 ? 2'h3 : io_n_in_9; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_en_r ? _GEN_0 : io_n_in_9; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_9(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_10 == 2'h2 ? 2'h3 : io_n_in_10; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_en_r ? _GEN_0 : io_n_in_10; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_10(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_11 == 2'h2 ? 2'h3 : io_n_in_11; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_en_r ? _GEN_0 : io_n_in_11; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_11(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_12 == 2'h2 ? 2'h3 : io_n_in_12; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_en_r ? _GEN_0 : io_n_in_12; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_12(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_13 == 2'h2 ? 2'h3 : io_n_in_13; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_en_r ? _GEN_0 : io_n_in_13; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_13(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_14 == 2'h2 ? 2'h3 : io_n_in_14; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_en_r ? _GEN_0 : io_n_in_14; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_14(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_15 == 2'h2 ? 2'h3 : io_n_in_15; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_en_r ? _GEN_0 : io_n_in_15; // @[router.scala 29:14 node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Exit_15(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_16 == 2'h2 ? 2'h3 : io_n_in_16; // @[router.scala 30:23 31:13 node.scala 30:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_en_r ? _GEN_0 : io_n_in_16; // @[router.scala 29:14 node.scala 30:9]
  assign io_x_out = io_x_in; // @[node.scala 31:9]
endmodule
module Idle(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_1 == 2'h3 ? 2'h0 : io_n_in_1; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_1 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_en_r ? _GEN_0 : io_n_in_1; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_1(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_2 == 2'h3 ? 2'h0 : io_n_in_2; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_2 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_en_r ? _GEN_0 : io_n_in_2; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_2(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_3 == 2'h3 ? 2'h0 : io_n_in_3; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_3 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_en_r ? _GEN_0 : io_n_in_3; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_3(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_4 == 2'h3 ? 2'h0 : io_n_in_4; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_4 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_en_r ? _GEN_0 : io_n_in_4; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_4(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_5 == 2'h3 ? 2'h0 : io_n_in_5; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_5 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_en_r ? _GEN_0 : io_n_in_5; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_5(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_6 == 2'h3 ? 2'h0 : io_n_in_6; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_6 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_en_r ? _GEN_0 : io_n_in_6; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_6(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_7 == 2'h3 ? 2'h0 : io_n_in_7; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_7 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_en_r ? _GEN_0 : io_n_in_7; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_7(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_8 == 2'h3 ? 2'h0 : io_n_in_8; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_8 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_en_r ? _GEN_0 : io_n_in_8; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_8(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_9 == 2'h3 ? 2'h0 : io_n_in_9; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_9 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_en_r ? _GEN_0 : io_n_in_9; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_9(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_10 == 2'h3 ? 2'h0 : io_n_in_10; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_10 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_en_r ? _GEN_0 : io_n_in_10; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_10(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_11 == 2'h3 ? 2'h0 : io_n_in_11; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_11 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_en_r ? _GEN_0 : io_n_in_11; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_11(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_12 == 2'h3 ? 2'h0 : io_n_in_12; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_12 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_en_r ? _GEN_0 : io_n_in_12; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_12(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_13 == 2'h3 ? 2'h0 : io_n_in_13; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_13 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_en_r ? _GEN_0 : io_n_in_13; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_13(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_14 == 2'h3 ? 2'h0 : io_n_in_14; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_14 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_en_r ? _GEN_0 : io_n_in_14; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_14(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_15 == 2'h3 ? 2'h0 : io_n_in_15; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_15 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_en_r ? _GEN_0 : io_n_in_15; // @[router.scala 36:14 node.scala 30:9]
  assign io_n_out_16 = io_n_in_16; // @[node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module Idle_15(
  input        io_en_r,
  input  [1:0] io_n_in_0,
  input  [1:0] io_n_in_1,
  input  [1:0] io_n_in_2,
  input  [1:0] io_n_in_3,
  input  [1:0] io_n_in_4,
  input  [1:0] io_n_in_5,
  input  [1:0] io_n_in_6,
  input  [1:0] io_n_in_7,
  input  [1:0] io_n_in_8,
  input  [1:0] io_n_in_9,
  input  [1:0] io_n_in_10,
  input  [1:0] io_n_in_11,
  input  [1:0] io_n_in_12,
  input  [1:0] io_n_in_13,
  input  [1:0] io_n_in_14,
  input  [1:0] io_n_in_15,
  input  [1:0] io_n_in_16,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  input        io_x_in,
  output       io_x_out
);
  wire [1:0] _GEN_0 = io_n_in_16 == 2'h3 ? 2'h0 : io_n_in_16; // @[router.scala 37:23 38:13 node.scala 30:9]
  wire  _GEN_1 = io_n_in_16 == 2'h3 | io_x_in; // @[router.scala 37:23 39:10 node.scala 31:9]
  assign io_n_out_0 = io_n_in_0; // @[node.scala 30:9]
  assign io_n_out_1 = io_n_in_1; // @[node.scala 30:9]
  assign io_n_out_2 = io_n_in_2; // @[node.scala 30:9]
  assign io_n_out_3 = io_n_in_3; // @[node.scala 30:9]
  assign io_n_out_4 = io_n_in_4; // @[node.scala 30:9]
  assign io_n_out_5 = io_n_in_5; // @[node.scala 30:9]
  assign io_n_out_6 = io_n_in_6; // @[node.scala 30:9]
  assign io_n_out_7 = io_n_in_7; // @[node.scala 30:9]
  assign io_n_out_8 = io_n_in_8; // @[node.scala 30:9]
  assign io_n_out_9 = io_n_in_9; // @[node.scala 30:9]
  assign io_n_out_10 = io_n_in_10; // @[node.scala 30:9]
  assign io_n_out_11 = io_n_in_11; // @[node.scala 30:9]
  assign io_n_out_12 = io_n_in_12; // @[node.scala 30:9]
  assign io_n_out_13 = io_n_in_13; // @[node.scala 30:9]
  assign io_n_out_14 = io_n_in_14; // @[node.scala 30:9]
  assign io_n_out_15 = io_n_in_15; // @[node.scala 30:9]
  assign io_n_out_16 = io_en_r ? _GEN_0 : io_n_in_16; // @[router.scala 36:14 node.scala 30:9]
  assign io_x_out = io_en_r ? _GEN_1 : io_x_in; // @[router.scala 36:14 node.scala 31:9]
endmodule
module system(
  input        clock,
  input        reset,
  input  [6:0] io_en_a,
  output [1:0] io_n_out_0,
  output [1:0] io_n_out_1,
  output [1:0] io_n_out_2,
  output [1:0] io_n_out_3,
  output [1:0] io_n_out_4,
  output [1:0] io_n_out_5,
  output [1:0] io_n_out_6,
  output [1:0] io_n_out_7,
  output [1:0] io_n_out_8,
  output [1:0] io_n_out_9,
  output [1:0] io_n_out_10,
  output [1:0] io_n_out_11,
  output [1:0] io_n_out_12,
  output [1:0] io_n_out_13,
  output [1:0] io_n_out_14,
  output [1:0] io_n_out_15,
  output [1:0] io_n_out_16,
  output       io_x_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rules_0_io_en_r; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_0; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_1; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_2; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_3; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_4; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_5; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_6; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_7; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_8; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_9; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_10; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_11; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_12; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_13; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_14; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_15; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_in_16; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_0; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_1; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_2; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_3; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_4; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_5; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_6; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_7; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_8; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_9; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_10; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_11; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_12; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_13; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_14; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_15; // @[system.scala 16:16]
  wire [1:0] rules_0_io_n_out_16; // @[system.scala 16:16]
  wire  rules_0_io_x_in; // @[system.scala 16:16]
  wire  rules_0_io_x_out; // @[system.scala 16:16]
  wire  rules_1_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_1_io_n_out_16; // @[system.scala 18:16]
  wire  rules_1_io_x_in; // @[system.scala 18:16]
  wire  rules_1_io_x_out; // @[system.scala 18:16]
  wire  rules_2_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_2_io_n_out_16; // @[system.scala 18:16]
  wire  rules_2_io_x_in; // @[system.scala 18:16]
  wire  rules_2_io_x_out; // @[system.scala 18:16]
  wire  rules_3_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_3_io_n_out_16; // @[system.scala 18:16]
  wire  rules_3_io_x_in; // @[system.scala 18:16]
  wire  rules_3_io_x_out; // @[system.scala 18:16]
  wire  rules_4_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_4_io_n_out_16; // @[system.scala 18:16]
  wire  rules_4_io_x_in; // @[system.scala 18:16]
  wire  rules_4_io_x_out; // @[system.scala 18:16]
  wire  rules_5_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_5_io_n_out_16; // @[system.scala 18:16]
  wire  rules_5_io_x_in; // @[system.scala 18:16]
  wire  rules_5_io_x_out; // @[system.scala 18:16]
  wire  rules_6_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_6_io_n_out_16; // @[system.scala 18:16]
  wire  rules_6_io_x_in; // @[system.scala 18:16]
  wire  rules_6_io_x_out; // @[system.scala 18:16]
  wire  rules_7_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_7_io_n_out_16; // @[system.scala 18:16]
  wire  rules_7_io_x_in; // @[system.scala 18:16]
  wire  rules_7_io_x_out; // @[system.scala 18:16]
  wire  rules_8_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_8_io_n_out_16; // @[system.scala 18:16]
  wire  rules_8_io_x_in; // @[system.scala 18:16]
  wire  rules_8_io_x_out; // @[system.scala 18:16]
  wire  rules_9_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_9_io_n_out_16; // @[system.scala 18:16]
  wire  rules_9_io_x_in; // @[system.scala 18:16]
  wire  rules_9_io_x_out; // @[system.scala 18:16]
  wire  rules_10_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_10_io_n_out_16; // @[system.scala 18:16]
  wire  rules_10_io_x_in; // @[system.scala 18:16]
  wire  rules_10_io_x_out; // @[system.scala 18:16]
  wire  rules_11_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_11_io_n_out_16; // @[system.scala 18:16]
  wire  rules_11_io_x_in; // @[system.scala 18:16]
  wire  rules_11_io_x_out; // @[system.scala 18:16]
  wire  rules_12_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_12_io_n_out_16; // @[system.scala 18:16]
  wire  rules_12_io_x_in; // @[system.scala 18:16]
  wire  rules_12_io_x_out; // @[system.scala 18:16]
  wire  rules_13_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_13_io_n_out_16; // @[system.scala 18:16]
  wire  rules_13_io_x_in; // @[system.scala 18:16]
  wire  rules_13_io_x_out; // @[system.scala 18:16]
  wire  rules_14_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_14_io_n_out_16; // @[system.scala 18:16]
  wire  rules_14_io_x_in; // @[system.scala 18:16]
  wire  rules_14_io_x_out; // @[system.scala 18:16]
  wire  rules_15_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_15_io_n_out_16; // @[system.scala 18:16]
  wire  rules_15_io_x_in; // @[system.scala 18:16]
  wire  rules_15_io_x_out; // @[system.scala 18:16]
  wire  rules_16_io_en_r; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_0; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_1; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_2; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_3; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_4; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_5; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_6; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_7; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_8; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_9; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_10; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_11; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_12; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_13; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_14; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_15; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_in_16; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_0; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_1; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_2; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_3; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_4; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_5; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_6; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_7; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_8; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_9; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_10; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_11; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_12; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_13; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_14; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_15; // @[system.scala 18:16]
  wire [1:0] rules_16_io_n_out_16; // @[system.scala 18:16]
  wire  rules_16_io_x_in; // @[system.scala 18:16]
  wire  rules_16_io_x_out; // @[system.scala 18:16]
  wire  rules_17_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_17_io_n_out_16; // @[system.scala 21:16]
  wire  rules_17_io_x_in; // @[system.scala 21:16]
  wire  rules_17_io_x_out; // @[system.scala 21:16]
  wire  rules_18_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_18_io_n_out_16; // @[system.scala 21:16]
  wire  rules_18_io_x_in; // @[system.scala 21:16]
  wire  rules_18_io_x_out; // @[system.scala 21:16]
  wire  rules_19_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_19_io_n_out_16; // @[system.scala 21:16]
  wire  rules_19_io_x_in; // @[system.scala 21:16]
  wire  rules_19_io_x_out; // @[system.scala 21:16]
  wire  rules_20_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_20_io_n_out_16; // @[system.scala 21:16]
  wire  rules_20_io_x_in; // @[system.scala 21:16]
  wire  rules_20_io_x_out; // @[system.scala 21:16]
  wire  rules_21_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_21_io_n_out_16; // @[system.scala 21:16]
  wire  rules_21_io_x_in; // @[system.scala 21:16]
  wire  rules_21_io_x_out; // @[system.scala 21:16]
  wire  rules_22_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_22_io_n_out_16; // @[system.scala 21:16]
  wire  rules_22_io_x_in; // @[system.scala 21:16]
  wire  rules_22_io_x_out; // @[system.scala 21:16]
  wire  rules_23_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_23_io_n_out_16; // @[system.scala 21:16]
  wire  rules_23_io_x_in; // @[system.scala 21:16]
  wire  rules_23_io_x_out; // @[system.scala 21:16]
  wire  rules_24_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_24_io_n_out_16; // @[system.scala 21:16]
  wire  rules_24_io_x_in; // @[system.scala 21:16]
  wire  rules_24_io_x_out; // @[system.scala 21:16]
  wire  rules_25_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_25_io_n_out_16; // @[system.scala 21:16]
  wire  rules_25_io_x_in; // @[system.scala 21:16]
  wire  rules_25_io_x_out; // @[system.scala 21:16]
  wire  rules_26_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_26_io_n_out_16; // @[system.scala 21:16]
  wire  rules_26_io_x_in; // @[system.scala 21:16]
  wire  rules_26_io_x_out; // @[system.scala 21:16]
  wire  rules_27_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_27_io_n_out_16; // @[system.scala 21:16]
  wire  rules_27_io_x_in; // @[system.scala 21:16]
  wire  rules_27_io_x_out; // @[system.scala 21:16]
  wire  rules_28_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_28_io_n_out_16; // @[system.scala 21:16]
  wire  rules_28_io_x_in; // @[system.scala 21:16]
  wire  rules_28_io_x_out; // @[system.scala 21:16]
  wire  rules_29_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_29_io_n_out_16; // @[system.scala 21:16]
  wire  rules_29_io_x_in; // @[system.scala 21:16]
  wire  rules_29_io_x_out; // @[system.scala 21:16]
  wire  rules_30_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_30_io_n_out_16; // @[system.scala 21:16]
  wire  rules_30_io_x_in; // @[system.scala 21:16]
  wire  rules_30_io_x_out; // @[system.scala 21:16]
  wire  rules_31_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_31_io_n_out_16; // @[system.scala 21:16]
  wire  rules_31_io_x_in; // @[system.scala 21:16]
  wire  rules_31_io_x_out; // @[system.scala 21:16]
  wire  rules_32_io_en_r; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_0; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_1; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_2; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_3; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_4; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_5; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_6; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_7; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_8; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_9; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_10; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_11; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_12; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_13; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_14; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_15; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_in_16; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_0; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_1; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_2; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_3; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_4; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_5; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_6; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_7; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_8; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_9; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_10; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_11; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_12; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_13; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_14; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_15; // @[system.scala 21:16]
  wire [1:0] rules_32_io_n_out_16; // @[system.scala 21:16]
  wire  rules_32_io_x_in; // @[system.scala 21:16]
  wire  rules_32_io_x_out; // @[system.scala 21:16]
  wire  rules_33_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_33_io_n_out_16; // @[system.scala 24:16]
  wire  rules_33_io_x_in; // @[system.scala 24:16]
  wire  rules_33_io_x_out; // @[system.scala 24:16]
  wire  rules_34_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_34_io_n_out_16; // @[system.scala 24:16]
  wire  rules_34_io_x_in; // @[system.scala 24:16]
  wire  rules_34_io_x_out; // @[system.scala 24:16]
  wire  rules_35_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_35_io_n_out_16; // @[system.scala 24:16]
  wire  rules_35_io_x_in; // @[system.scala 24:16]
  wire  rules_35_io_x_out; // @[system.scala 24:16]
  wire  rules_36_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_36_io_n_out_16; // @[system.scala 24:16]
  wire  rules_36_io_x_in; // @[system.scala 24:16]
  wire  rules_36_io_x_out; // @[system.scala 24:16]
  wire  rules_37_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_37_io_n_out_16; // @[system.scala 24:16]
  wire  rules_37_io_x_in; // @[system.scala 24:16]
  wire  rules_37_io_x_out; // @[system.scala 24:16]
  wire  rules_38_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_38_io_n_out_16; // @[system.scala 24:16]
  wire  rules_38_io_x_in; // @[system.scala 24:16]
  wire  rules_38_io_x_out; // @[system.scala 24:16]
  wire  rules_39_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_39_io_n_out_16; // @[system.scala 24:16]
  wire  rules_39_io_x_in; // @[system.scala 24:16]
  wire  rules_39_io_x_out; // @[system.scala 24:16]
  wire  rules_40_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_40_io_n_out_16; // @[system.scala 24:16]
  wire  rules_40_io_x_in; // @[system.scala 24:16]
  wire  rules_40_io_x_out; // @[system.scala 24:16]
  wire  rules_41_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_41_io_n_out_16; // @[system.scala 24:16]
  wire  rules_41_io_x_in; // @[system.scala 24:16]
  wire  rules_41_io_x_out; // @[system.scala 24:16]
  wire  rules_42_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_42_io_n_out_16; // @[system.scala 24:16]
  wire  rules_42_io_x_in; // @[system.scala 24:16]
  wire  rules_42_io_x_out; // @[system.scala 24:16]
  wire  rules_43_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_43_io_n_out_16; // @[system.scala 24:16]
  wire  rules_43_io_x_in; // @[system.scala 24:16]
  wire  rules_43_io_x_out; // @[system.scala 24:16]
  wire  rules_44_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_44_io_n_out_16; // @[system.scala 24:16]
  wire  rules_44_io_x_in; // @[system.scala 24:16]
  wire  rules_44_io_x_out; // @[system.scala 24:16]
  wire  rules_45_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_45_io_n_out_16; // @[system.scala 24:16]
  wire  rules_45_io_x_in; // @[system.scala 24:16]
  wire  rules_45_io_x_out; // @[system.scala 24:16]
  wire  rules_46_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_46_io_n_out_16; // @[system.scala 24:16]
  wire  rules_46_io_x_in; // @[system.scala 24:16]
  wire  rules_46_io_x_out; // @[system.scala 24:16]
  wire  rules_47_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_47_io_n_out_16; // @[system.scala 24:16]
  wire  rules_47_io_x_in; // @[system.scala 24:16]
  wire  rules_47_io_x_out; // @[system.scala 24:16]
  wire  rules_48_io_en_r; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_0; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_1; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_2; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_3; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_4; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_5; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_6; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_7; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_8; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_9; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_10; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_11; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_12; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_13; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_14; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_15; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_in_16; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_0; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_1; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_2; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_3; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_4; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_5; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_6; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_7; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_8; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_9; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_10; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_11; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_12; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_13; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_14; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_15; // @[system.scala 24:16]
  wire [1:0] rules_48_io_n_out_16; // @[system.scala 24:16]
  wire  rules_48_io_x_in; // @[system.scala 24:16]
  wire  rules_48_io_x_out; // @[system.scala 24:16]
  wire  rules_49_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_49_io_n_out_16; // @[system.scala 27:16]
  wire  rules_49_io_x_in; // @[system.scala 27:16]
  wire  rules_49_io_x_out; // @[system.scala 27:16]
  wire  rules_50_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_50_io_n_out_16; // @[system.scala 27:16]
  wire  rules_50_io_x_in; // @[system.scala 27:16]
  wire  rules_50_io_x_out; // @[system.scala 27:16]
  wire  rules_51_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_51_io_n_out_16; // @[system.scala 27:16]
  wire  rules_51_io_x_in; // @[system.scala 27:16]
  wire  rules_51_io_x_out; // @[system.scala 27:16]
  wire  rules_52_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_52_io_n_out_16; // @[system.scala 27:16]
  wire  rules_52_io_x_in; // @[system.scala 27:16]
  wire  rules_52_io_x_out; // @[system.scala 27:16]
  wire  rules_53_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_53_io_n_out_16; // @[system.scala 27:16]
  wire  rules_53_io_x_in; // @[system.scala 27:16]
  wire  rules_53_io_x_out; // @[system.scala 27:16]
  wire  rules_54_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_54_io_n_out_16; // @[system.scala 27:16]
  wire  rules_54_io_x_in; // @[system.scala 27:16]
  wire  rules_54_io_x_out; // @[system.scala 27:16]
  wire  rules_55_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_55_io_n_out_16; // @[system.scala 27:16]
  wire  rules_55_io_x_in; // @[system.scala 27:16]
  wire  rules_55_io_x_out; // @[system.scala 27:16]
  wire  rules_56_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_56_io_n_out_16; // @[system.scala 27:16]
  wire  rules_56_io_x_in; // @[system.scala 27:16]
  wire  rules_56_io_x_out; // @[system.scala 27:16]
  wire  rules_57_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_57_io_n_out_16; // @[system.scala 27:16]
  wire  rules_57_io_x_in; // @[system.scala 27:16]
  wire  rules_57_io_x_out; // @[system.scala 27:16]
  wire  rules_58_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_58_io_n_out_16; // @[system.scala 27:16]
  wire  rules_58_io_x_in; // @[system.scala 27:16]
  wire  rules_58_io_x_out; // @[system.scala 27:16]
  wire  rules_59_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_59_io_n_out_16; // @[system.scala 27:16]
  wire  rules_59_io_x_in; // @[system.scala 27:16]
  wire  rules_59_io_x_out; // @[system.scala 27:16]
  wire  rules_60_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_60_io_n_out_16; // @[system.scala 27:16]
  wire  rules_60_io_x_in; // @[system.scala 27:16]
  wire  rules_60_io_x_out; // @[system.scala 27:16]
  wire  rules_61_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_61_io_n_out_16; // @[system.scala 27:16]
  wire  rules_61_io_x_in; // @[system.scala 27:16]
  wire  rules_61_io_x_out; // @[system.scala 27:16]
  wire  rules_62_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_62_io_n_out_16; // @[system.scala 27:16]
  wire  rules_62_io_x_in; // @[system.scala 27:16]
  wire  rules_62_io_x_out; // @[system.scala 27:16]
  wire  rules_63_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_63_io_n_out_16; // @[system.scala 27:16]
  wire  rules_63_io_x_in; // @[system.scala 27:16]
  wire  rules_63_io_x_out; // @[system.scala 27:16]
  wire  rules_64_io_en_r; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_0; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_1; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_2; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_3; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_4; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_5; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_6; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_7; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_8; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_9; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_10; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_11; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_12; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_13; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_14; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_15; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_in_16; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_0; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_1; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_2; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_3; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_4; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_5; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_6; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_7; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_8; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_9; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_10; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_11; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_12; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_13; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_14; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_15; // @[system.scala 27:16]
  wire [1:0] rules_64_io_n_out_16; // @[system.scala 27:16]
  wire  rules_64_io_x_in; // @[system.scala 27:16]
  wire  rules_64_io_x_out; // @[system.scala 27:16]
  reg [1:0] n_reg_0; // @[system.scala 12:16]
  reg [1:0] n_reg_1; // @[system.scala 12:16]
  reg [1:0] n_reg_2; // @[system.scala 12:16]
  reg [1:0] n_reg_3; // @[system.scala 12:16]
  reg [1:0] n_reg_4; // @[system.scala 12:16]
  reg [1:0] n_reg_5; // @[system.scala 12:16]
  reg [1:0] n_reg_6; // @[system.scala 12:16]
  reg [1:0] n_reg_7; // @[system.scala 12:16]
  reg [1:0] n_reg_8; // @[system.scala 12:16]
  reg [1:0] n_reg_9; // @[system.scala 12:16]
  reg [1:0] n_reg_10; // @[system.scala 12:16]
  reg [1:0] n_reg_11; // @[system.scala 12:16]
  reg [1:0] n_reg_12; // @[system.scala 12:16]
  reg [1:0] n_reg_13; // @[system.scala 12:16]
  reg [1:0] n_reg_14; // @[system.scala 12:16]
  reg [1:0] n_reg_15; // @[system.scala 12:16]
  reg [1:0] n_reg_16; // @[system.scala 12:16]
  reg  x_reg; // @[system.scala 14:16]
  wire  _T = io_en_a == 7'h0; // @[system.scala 32:27]
  wire [1:0] _GEN_0 = _T ? rules_0_io_n_out_0 : n_reg_0; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_1 = _T ? rules_0_io_n_out_1 : n_reg_1; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_2 = _T ? rules_0_io_n_out_2 : n_reg_2; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_3 = _T ? rules_0_io_n_out_3 : n_reg_3; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_4 = _T ? rules_0_io_n_out_4 : n_reg_4; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_5 = _T ? rules_0_io_n_out_5 : n_reg_5; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_6 = _T ? rules_0_io_n_out_6 : n_reg_6; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_7 = _T ? rules_0_io_n_out_7 : n_reg_7; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_8 = _T ? rules_0_io_n_out_8 : n_reg_8; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_9 = _T ? rules_0_io_n_out_9 : n_reg_9; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_10 = _T ? rules_0_io_n_out_10 : n_reg_10; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_11 = _T ? rules_0_io_n_out_11 : n_reg_11; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_12 = _T ? rules_0_io_n_out_12 : n_reg_12; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_13 = _T ? rules_0_io_n_out_13 : n_reg_13; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_14 = _T ? rules_0_io_n_out_14 : n_reg_14; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_15 = _T ? rules_0_io_n_out_15 : n_reg_15; // @[system.scala 12:16 33:21 34:7]
  wire [1:0] _GEN_16 = _T ? rules_0_io_n_out_16 : n_reg_16; // @[system.scala 12:16 33:21 34:7]
  wire  _GEN_17 = _T ? rules_0_io_x_out : x_reg; // @[system.scala 14:16 33:21 35:7]
  wire  _T_2 = io_en_a == 7'h1; // @[system.scala 32:27]
  wire [1:0] _GEN_18 = _T_2 ? rules_1_io_n_out_0 : _GEN_0; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_19 = _T_2 ? rules_1_io_n_out_1 : _GEN_1; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_20 = _T_2 ? rules_1_io_n_out_2 : _GEN_2; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_21 = _T_2 ? rules_1_io_n_out_3 : _GEN_3; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_22 = _T_2 ? rules_1_io_n_out_4 : _GEN_4; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_23 = _T_2 ? rules_1_io_n_out_5 : _GEN_5; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_24 = _T_2 ? rules_1_io_n_out_6 : _GEN_6; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_25 = _T_2 ? rules_1_io_n_out_7 : _GEN_7; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_26 = _T_2 ? rules_1_io_n_out_8 : _GEN_8; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_27 = _T_2 ? rules_1_io_n_out_9 : _GEN_9; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_28 = _T_2 ? rules_1_io_n_out_10 : _GEN_10; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_29 = _T_2 ? rules_1_io_n_out_11 : _GEN_11; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_30 = _T_2 ? rules_1_io_n_out_12 : _GEN_12; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_31 = _T_2 ? rules_1_io_n_out_13 : _GEN_13; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_32 = _T_2 ? rules_1_io_n_out_14 : _GEN_14; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_33 = _T_2 ? rules_1_io_n_out_15 : _GEN_15; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_34 = _T_2 ? rules_1_io_n_out_16 : _GEN_16; // @[system.scala 33:21 34:7]
  wire  _GEN_35 = _T_2 ? rules_1_io_x_out : _GEN_17; // @[system.scala 33:21 35:7]
  wire  _T_4 = io_en_a == 7'h2; // @[system.scala 32:27]
  wire [1:0] _GEN_36 = _T_4 ? rules_2_io_n_out_0 : _GEN_18; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_37 = _T_4 ? rules_2_io_n_out_1 : _GEN_19; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_38 = _T_4 ? rules_2_io_n_out_2 : _GEN_20; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_39 = _T_4 ? rules_2_io_n_out_3 : _GEN_21; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_40 = _T_4 ? rules_2_io_n_out_4 : _GEN_22; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_41 = _T_4 ? rules_2_io_n_out_5 : _GEN_23; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_42 = _T_4 ? rules_2_io_n_out_6 : _GEN_24; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_43 = _T_4 ? rules_2_io_n_out_7 : _GEN_25; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_44 = _T_4 ? rules_2_io_n_out_8 : _GEN_26; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_45 = _T_4 ? rules_2_io_n_out_9 : _GEN_27; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_46 = _T_4 ? rules_2_io_n_out_10 : _GEN_28; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_47 = _T_4 ? rules_2_io_n_out_11 : _GEN_29; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_48 = _T_4 ? rules_2_io_n_out_12 : _GEN_30; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_49 = _T_4 ? rules_2_io_n_out_13 : _GEN_31; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_50 = _T_4 ? rules_2_io_n_out_14 : _GEN_32; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_51 = _T_4 ? rules_2_io_n_out_15 : _GEN_33; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_52 = _T_4 ? rules_2_io_n_out_16 : _GEN_34; // @[system.scala 33:21 34:7]
  wire  _GEN_53 = _T_4 ? rules_2_io_x_out : _GEN_35; // @[system.scala 33:21 35:7]
  wire  _T_6 = io_en_a == 7'h3; // @[system.scala 32:27]
  wire [1:0] _GEN_54 = _T_6 ? rules_3_io_n_out_0 : _GEN_36; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_55 = _T_6 ? rules_3_io_n_out_1 : _GEN_37; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_56 = _T_6 ? rules_3_io_n_out_2 : _GEN_38; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_57 = _T_6 ? rules_3_io_n_out_3 : _GEN_39; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_58 = _T_6 ? rules_3_io_n_out_4 : _GEN_40; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_59 = _T_6 ? rules_3_io_n_out_5 : _GEN_41; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_60 = _T_6 ? rules_3_io_n_out_6 : _GEN_42; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_61 = _T_6 ? rules_3_io_n_out_7 : _GEN_43; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_62 = _T_6 ? rules_3_io_n_out_8 : _GEN_44; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_63 = _T_6 ? rules_3_io_n_out_9 : _GEN_45; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_64 = _T_6 ? rules_3_io_n_out_10 : _GEN_46; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_65 = _T_6 ? rules_3_io_n_out_11 : _GEN_47; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_66 = _T_6 ? rules_3_io_n_out_12 : _GEN_48; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_67 = _T_6 ? rules_3_io_n_out_13 : _GEN_49; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_68 = _T_6 ? rules_3_io_n_out_14 : _GEN_50; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_69 = _T_6 ? rules_3_io_n_out_15 : _GEN_51; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_70 = _T_6 ? rules_3_io_n_out_16 : _GEN_52; // @[system.scala 33:21 34:7]
  wire  _GEN_71 = _T_6 ? rules_3_io_x_out : _GEN_53; // @[system.scala 33:21 35:7]
  wire  _T_8 = io_en_a == 7'h4; // @[system.scala 32:27]
  wire [1:0] _GEN_72 = _T_8 ? rules_4_io_n_out_0 : _GEN_54; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_73 = _T_8 ? rules_4_io_n_out_1 : _GEN_55; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_74 = _T_8 ? rules_4_io_n_out_2 : _GEN_56; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_75 = _T_8 ? rules_4_io_n_out_3 : _GEN_57; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_76 = _T_8 ? rules_4_io_n_out_4 : _GEN_58; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_77 = _T_8 ? rules_4_io_n_out_5 : _GEN_59; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_78 = _T_8 ? rules_4_io_n_out_6 : _GEN_60; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_79 = _T_8 ? rules_4_io_n_out_7 : _GEN_61; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_80 = _T_8 ? rules_4_io_n_out_8 : _GEN_62; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_81 = _T_8 ? rules_4_io_n_out_9 : _GEN_63; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_82 = _T_8 ? rules_4_io_n_out_10 : _GEN_64; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_83 = _T_8 ? rules_4_io_n_out_11 : _GEN_65; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_84 = _T_8 ? rules_4_io_n_out_12 : _GEN_66; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_85 = _T_8 ? rules_4_io_n_out_13 : _GEN_67; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_86 = _T_8 ? rules_4_io_n_out_14 : _GEN_68; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_87 = _T_8 ? rules_4_io_n_out_15 : _GEN_69; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_88 = _T_8 ? rules_4_io_n_out_16 : _GEN_70; // @[system.scala 33:21 34:7]
  wire  _GEN_89 = _T_8 ? rules_4_io_x_out : _GEN_71; // @[system.scala 33:21 35:7]
  wire  _T_10 = io_en_a == 7'h5; // @[system.scala 32:27]
  wire [1:0] _GEN_90 = _T_10 ? rules_5_io_n_out_0 : _GEN_72; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_91 = _T_10 ? rules_5_io_n_out_1 : _GEN_73; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_92 = _T_10 ? rules_5_io_n_out_2 : _GEN_74; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_93 = _T_10 ? rules_5_io_n_out_3 : _GEN_75; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_94 = _T_10 ? rules_5_io_n_out_4 : _GEN_76; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_95 = _T_10 ? rules_5_io_n_out_5 : _GEN_77; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_96 = _T_10 ? rules_5_io_n_out_6 : _GEN_78; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_97 = _T_10 ? rules_5_io_n_out_7 : _GEN_79; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_98 = _T_10 ? rules_5_io_n_out_8 : _GEN_80; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_99 = _T_10 ? rules_5_io_n_out_9 : _GEN_81; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_100 = _T_10 ? rules_5_io_n_out_10 : _GEN_82; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_101 = _T_10 ? rules_5_io_n_out_11 : _GEN_83; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_102 = _T_10 ? rules_5_io_n_out_12 : _GEN_84; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_103 = _T_10 ? rules_5_io_n_out_13 : _GEN_85; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_104 = _T_10 ? rules_5_io_n_out_14 : _GEN_86; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_105 = _T_10 ? rules_5_io_n_out_15 : _GEN_87; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_106 = _T_10 ? rules_5_io_n_out_16 : _GEN_88; // @[system.scala 33:21 34:7]
  wire  _GEN_107 = _T_10 ? rules_5_io_x_out : _GEN_89; // @[system.scala 33:21 35:7]
  wire  _T_12 = io_en_a == 7'h6; // @[system.scala 32:27]
  wire [1:0] _GEN_108 = _T_12 ? rules_6_io_n_out_0 : _GEN_90; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_109 = _T_12 ? rules_6_io_n_out_1 : _GEN_91; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_110 = _T_12 ? rules_6_io_n_out_2 : _GEN_92; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_111 = _T_12 ? rules_6_io_n_out_3 : _GEN_93; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_112 = _T_12 ? rules_6_io_n_out_4 : _GEN_94; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_113 = _T_12 ? rules_6_io_n_out_5 : _GEN_95; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_114 = _T_12 ? rules_6_io_n_out_6 : _GEN_96; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_115 = _T_12 ? rules_6_io_n_out_7 : _GEN_97; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_116 = _T_12 ? rules_6_io_n_out_8 : _GEN_98; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_117 = _T_12 ? rules_6_io_n_out_9 : _GEN_99; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_118 = _T_12 ? rules_6_io_n_out_10 : _GEN_100; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_119 = _T_12 ? rules_6_io_n_out_11 : _GEN_101; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_120 = _T_12 ? rules_6_io_n_out_12 : _GEN_102; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_121 = _T_12 ? rules_6_io_n_out_13 : _GEN_103; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_122 = _T_12 ? rules_6_io_n_out_14 : _GEN_104; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_123 = _T_12 ? rules_6_io_n_out_15 : _GEN_105; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_124 = _T_12 ? rules_6_io_n_out_16 : _GEN_106; // @[system.scala 33:21 34:7]
  wire  _GEN_125 = _T_12 ? rules_6_io_x_out : _GEN_107; // @[system.scala 33:21 35:7]
  wire  _T_14 = io_en_a == 7'h7; // @[system.scala 32:27]
  wire [1:0] _GEN_126 = _T_14 ? rules_7_io_n_out_0 : _GEN_108; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_127 = _T_14 ? rules_7_io_n_out_1 : _GEN_109; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_128 = _T_14 ? rules_7_io_n_out_2 : _GEN_110; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_129 = _T_14 ? rules_7_io_n_out_3 : _GEN_111; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_130 = _T_14 ? rules_7_io_n_out_4 : _GEN_112; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_131 = _T_14 ? rules_7_io_n_out_5 : _GEN_113; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_132 = _T_14 ? rules_7_io_n_out_6 : _GEN_114; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_133 = _T_14 ? rules_7_io_n_out_7 : _GEN_115; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_134 = _T_14 ? rules_7_io_n_out_8 : _GEN_116; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_135 = _T_14 ? rules_7_io_n_out_9 : _GEN_117; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_136 = _T_14 ? rules_7_io_n_out_10 : _GEN_118; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_137 = _T_14 ? rules_7_io_n_out_11 : _GEN_119; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_138 = _T_14 ? rules_7_io_n_out_12 : _GEN_120; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_139 = _T_14 ? rules_7_io_n_out_13 : _GEN_121; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_140 = _T_14 ? rules_7_io_n_out_14 : _GEN_122; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_141 = _T_14 ? rules_7_io_n_out_15 : _GEN_123; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_142 = _T_14 ? rules_7_io_n_out_16 : _GEN_124; // @[system.scala 33:21 34:7]
  wire  _GEN_143 = _T_14 ? rules_7_io_x_out : _GEN_125; // @[system.scala 33:21 35:7]
  wire  _T_16 = io_en_a == 7'h8; // @[system.scala 32:27]
  wire [1:0] _GEN_144 = _T_16 ? rules_8_io_n_out_0 : _GEN_126; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_145 = _T_16 ? rules_8_io_n_out_1 : _GEN_127; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_146 = _T_16 ? rules_8_io_n_out_2 : _GEN_128; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_147 = _T_16 ? rules_8_io_n_out_3 : _GEN_129; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_148 = _T_16 ? rules_8_io_n_out_4 : _GEN_130; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_149 = _T_16 ? rules_8_io_n_out_5 : _GEN_131; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_150 = _T_16 ? rules_8_io_n_out_6 : _GEN_132; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_151 = _T_16 ? rules_8_io_n_out_7 : _GEN_133; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_152 = _T_16 ? rules_8_io_n_out_8 : _GEN_134; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_153 = _T_16 ? rules_8_io_n_out_9 : _GEN_135; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_154 = _T_16 ? rules_8_io_n_out_10 : _GEN_136; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_155 = _T_16 ? rules_8_io_n_out_11 : _GEN_137; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_156 = _T_16 ? rules_8_io_n_out_12 : _GEN_138; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_157 = _T_16 ? rules_8_io_n_out_13 : _GEN_139; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_158 = _T_16 ? rules_8_io_n_out_14 : _GEN_140; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_159 = _T_16 ? rules_8_io_n_out_15 : _GEN_141; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_160 = _T_16 ? rules_8_io_n_out_16 : _GEN_142; // @[system.scala 33:21 34:7]
  wire  _GEN_161 = _T_16 ? rules_8_io_x_out : _GEN_143; // @[system.scala 33:21 35:7]
  wire  _T_18 = io_en_a == 7'h9; // @[system.scala 32:27]
  wire [1:0] _GEN_162 = _T_18 ? rules_9_io_n_out_0 : _GEN_144; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_163 = _T_18 ? rules_9_io_n_out_1 : _GEN_145; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_164 = _T_18 ? rules_9_io_n_out_2 : _GEN_146; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_165 = _T_18 ? rules_9_io_n_out_3 : _GEN_147; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_166 = _T_18 ? rules_9_io_n_out_4 : _GEN_148; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_167 = _T_18 ? rules_9_io_n_out_5 : _GEN_149; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_168 = _T_18 ? rules_9_io_n_out_6 : _GEN_150; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_169 = _T_18 ? rules_9_io_n_out_7 : _GEN_151; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_170 = _T_18 ? rules_9_io_n_out_8 : _GEN_152; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_171 = _T_18 ? rules_9_io_n_out_9 : _GEN_153; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_172 = _T_18 ? rules_9_io_n_out_10 : _GEN_154; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_173 = _T_18 ? rules_9_io_n_out_11 : _GEN_155; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_174 = _T_18 ? rules_9_io_n_out_12 : _GEN_156; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_175 = _T_18 ? rules_9_io_n_out_13 : _GEN_157; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_176 = _T_18 ? rules_9_io_n_out_14 : _GEN_158; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_177 = _T_18 ? rules_9_io_n_out_15 : _GEN_159; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_178 = _T_18 ? rules_9_io_n_out_16 : _GEN_160; // @[system.scala 33:21 34:7]
  wire  _GEN_179 = _T_18 ? rules_9_io_x_out : _GEN_161; // @[system.scala 33:21 35:7]
  wire  _T_20 = io_en_a == 7'ha; // @[system.scala 32:27]
  wire [1:0] _GEN_180 = _T_20 ? rules_10_io_n_out_0 : _GEN_162; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_181 = _T_20 ? rules_10_io_n_out_1 : _GEN_163; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_182 = _T_20 ? rules_10_io_n_out_2 : _GEN_164; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_183 = _T_20 ? rules_10_io_n_out_3 : _GEN_165; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_184 = _T_20 ? rules_10_io_n_out_4 : _GEN_166; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_185 = _T_20 ? rules_10_io_n_out_5 : _GEN_167; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_186 = _T_20 ? rules_10_io_n_out_6 : _GEN_168; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_187 = _T_20 ? rules_10_io_n_out_7 : _GEN_169; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_188 = _T_20 ? rules_10_io_n_out_8 : _GEN_170; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_189 = _T_20 ? rules_10_io_n_out_9 : _GEN_171; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_190 = _T_20 ? rules_10_io_n_out_10 : _GEN_172; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_191 = _T_20 ? rules_10_io_n_out_11 : _GEN_173; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_192 = _T_20 ? rules_10_io_n_out_12 : _GEN_174; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_193 = _T_20 ? rules_10_io_n_out_13 : _GEN_175; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_194 = _T_20 ? rules_10_io_n_out_14 : _GEN_176; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_195 = _T_20 ? rules_10_io_n_out_15 : _GEN_177; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_196 = _T_20 ? rules_10_io_n_out_16 : _GEN_178; // @[system.scala 33:21 34:7]
  wire  _GEN_197 = _T_20 ? rules_10_io_x_out : _GEN_179; // @[system.scala 33:21 35:7]
  wire  _T_22 = io_en_a == 7'hb; // @[system.scala 32:27]
  wire [1:0] _GEN_198 = _T_22 ? rules_11_io_n_out_0 : _GEN_180; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_199 = _T_22 ? rules_11_io_n_out_1 : _GEN_181; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_200 = _T_22 ? rules_11_io_n_out_2 : _GEN_182; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_201 = _T_22 ? rules_11_io_n_out_3 : _GEN_183; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_202 = _T_22 ? rules_11_io_n_out_4 : _GEN_184; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_203 = _T_22 ? rules_11_io_n_out_5 : _GEN_185; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_204 = _T_22 ? rules_11_io_n_out_6 : _GEN_186; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_205 = _T_22 ? rules_11_io_n_out_7 : _GEN_187; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_206 = _T_22 ? rules_11_io_n_out_8 : _GEN_188; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_207 = _T_22 ? rules_11_io_n_out_9 : _GEN_189; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_208 = _T_22 ? rules_11_io_n_out_10 : _GEN_190; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_209 = _T_22 ? rules_11_io_n_out_11 : _GEN_191; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_210 = _T_22 ? rules_11_io_n_out_12 : _GEN_192; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_211 = _T_22 ? rules_11_io_n_out_13 : _GEN_193; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_212 = _T_22 ? rules_11_io_n_out_14 : _GEN_194; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_213 = _T_22 ? rules_11_io_n_out_15 : _GEN_195; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_214 = _T_22 ? rules_11_io_n_out_16 : _GEN_196; // @[system.scala 33:21 34:7]
  wire  _GEN_215 = _T_22 ? rules_11_io_x_out : _GEN_197; // @[system.scala 33:21 35:7]
  wire  _T_24 = io_en_a == 7'hc; // @[system.scala 32:27]
  wire [1:0] _GEN_216 = _T_24 ? rules_12_io_n_out_0 : _GEN_198; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_217 = _T_24 ? rules_12_io_n_out_1 : _GEN_199; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_218 = _T_24 ? rules_12_io_n_out_2 : _GEN_200; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_219 = _T_24 ? rules_12_io_n_out_3 : _GEN_201; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_220 = _T_24 ? rules_12_io_n_out_4 : _GEN_202; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_221 = _T_24 ? rules_12_io_n_out_5 : _GEN_203; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_222 = _T_24 ? rules_12_io_n_out_6 : _GEN_204; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_223 = _T_24 ? rules_12_io_n_out_7 : _GEN_205; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_224 = _T_24 ? rules_12_io_n_out_8 : _GEN_206; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_225 = _T_24 ? rules_12_io_n_out_9 : _GEN_207; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_226 = _T_24 ? rules_12_io_n_out_10 : _GEN_208; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_227 = _T_24 ? rules_12_io_n_out_11 : _GEN_209; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_228 = _T_24 ? rules_12_io_n_out_12 : _GEN_210; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_229 = _T_24 ? rules_12_io_n_out_13 : _GEN_211; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_230 = _T_24 ? rules_12_io_n_out_14 : _GEN_212; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_231 = _T_24 ? rules_12_io_n_out_15 : _GEN_213; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_232 = _T_24 ? rules_12_io_n_out_16 : _GEN_214; // @[system.scala 33:21 34:7]
  wire  _GEN_233 = _T_24 ? rules_12_io_x_out : _GEN_215; // @[system.scala 33:21 35:7]
  wire  _T_26 = io_en_a == 7'hd; // @[system.scala 32:27]
  wire [1:0] _GEN_234 = _T_26 ? rules_13_io_n_out_0 : _GEN_216; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_235 = _T_26 ? rules_13_io_n_out_1 : _GEN_217; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_236 = _T_26 ? rules_13_io_n_out_2 : _GEN_218; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_237 = _T_26 ? rules_13_io_n_out_3 : _GEN_219; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_238 = _T_26 ? rules_13_io_n_out_4 : _GEN_220; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_239 = _T_26 ? rules_13_io_n_out_5 : _GEN_221; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_240 = _T_26 ? rules_13_io_n_out_6 : _GEN_222; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_241 = _T_26 ? rules_13_io_n_out_7 : _GEN_223; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_242 = _T_26 ? rules_13_io_n_out_8 : _GEN_224; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_243 = _T_26 ? rules_13_io_n_out_9 : _GEN_225; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_244 = _T_26 ? rules_13_io_n_out_10 : _GEN_226; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_245 = _T_26 ? rules_13_io_n_out_11 : _GEN_227; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_246 = _T_26 ? rules_13_io_n_out_12 : _GEN_228; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_247 = _T_26 ? rules_13_io_n_out_13 : _GEN_229; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_248 = _T_26 ? rules_13_io_n_out_14 : _GEN_230; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_249 = _T_26 ? rules_13_io_n_out_15 : _GEN_231; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_250 = _T_26 ? rules_13_io_n_out_16 : _GEN_232; // @[system.scala 33:21 34:7]
  wire  _GEN_251 = _T_26 ? rules_13_io_x_out : _GEN_233; // @[system.scala 33:21 35:7]
  wire  _T_28 = io_en_a == 7'he; // @[system.scala 32:27]
  wire [1:0] _GEN_252 = _T_28 ? rules_14_io_n_out_0 : _GEN_234; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_253 = _T_28 ? rules_14_io_n_out_1 : _GEN_235; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_254 = _T_28 ? rules_14_io_n_out_2 : _GEN_236; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_255 = _T_28 ? rules_14_io_n_out_3 : _GEN_237; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_256 = _T_28 ? rules_14_io_n_out_4 : _GEN_238; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_257 = _T_28 ? rules_14_io_n_out_5 : _GEN_239; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_258 = _T_28 ? rules_14_io_n_out_6 : _GEN_240; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_259 = _T_28 ? rules_14_io_n_out_7 : _GEN_241; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_260 = _T_28 ? rules_14_io_n_out_8 : _GEN_242; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_261 = _T_28 ? rules_14_io_n_out_9 : _GEN_243; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_262 = _T_28 ? rules_14_io_n_out_10 : _GEN_244; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_263 = _T_28 ? rules_14_io_n_out_11 : _GEN_245; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_264 = _T_28 ? rules_14_io_n_out_12 : _GEN_246; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_265 = _T_28 ? rules_14_io_n_out_13 : _GEN_247; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_266 = _T_28 ? rules_14_io_n_out_14 : _GEN_248; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_267 = _T_28 ? rules_14_io_n_out_15 : _GEN_249; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_268 = _T_28 ? rules_14_io_n_out_16 : _GEN_250; // @[system.scala 33:21 34:7]
  wire  _GEN_269 = _T_28 ? rules_14_io_x_out : _GEN_251; // @[system.scala 33:21 35:7]
  wire  _T_30 = io_en_a == 7'hf; // @[system.scala 32:27]
  wire [1:0] _GEN_270 = _T_30 ? rules_15_io_n_out_0 : _GEN_252; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_271 = _T_30 ? rules_15_io_n_out_1 : _GEN_253; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_272 = _T_30 ? rules_15_io_n_out_2 : _GEN_254; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_273 = _T_30 ? rules_15_io_n_out_3 : _GEN_255; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_274 = _T_30 ? rules_15_io_n_out_4 : _GEN_256; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_275 = _T_30 ? rules_15_io_n_out_5 : _GEN_257; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_276 = _T_30 ? rules_15_io_n_out_6 : _GEN_258; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_277 = _T_30 ? rules_15_io_n_out_7 : _GEN_259; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_278 = _T_30 ? rules_15_io_n_out_8 : _GEN_260; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_279 = _T_30 ? rules_15_io_n_out_9 : _GEN_261; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_280 = _T_30 ? rules_15_io_n_out_10 : _GEN_262; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_281 = _T_30 ? rules_15_io_n_out_11 : _GEN_263; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_282 = _T_30 ? rules_15_io_n_out_12 : _GEN_264; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_283 = _T_30 ? rules_15_io_n_out_13 : _GEN_265; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_284 = _T_30 ? rules_15_io_n_out_14 : _GEN_266; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_285 = _T_30 ? rules_15_io_n_out_15 : _GEN_267; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_286 = _T_30 ? rules_15_io_n_out_16 : _GEN_268; // @[system.scala 33:21 34:7]
  wire  _GEN_287 = _T_30 ? rules_15_io_x_out : _GEN_269; // @[system.scala 33:21 35:7]
  wire  _T_32 = io_en_a == 7'h10; // @[system.scala 32:27]
  wire [1:0] _GEN_288 = _T_32 ? rules_16_io_n_out_0 : _GEN_270; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_289 = _T_32 ? rules_16_io_n_out_1 : _GEN_271; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_290 = _T_32 ? rules_16_io_n_out_2 : _GEN_272; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_291 = _T_32 ? rules_16_io_n_out_3 : _GEN_273; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_292 = _T_32 ? rules_16_io_n_out_4 : _GEN_274; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_293 = _T_32 ? rules_16_io_n_out_5 : _GEN_275; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_294 = _T_32 ? rules_16_io_n_out_6 : _GEN_276; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_295 = _T_32 ? rules_16_io_n_out_7 : _GEN_277; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_296 = _T_32 ? rules_16_io_n_out_8 : _GEN_278; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_297 = _T_32 ? rules_16_io_n_out_9 : _GEN_279; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_298 = _T_32 ? rules_16_io_n_out_10 : _GEN_280; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_299 = _T_32 ? rules_16_io_n_out_11 : _GEN_281; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_300 = _T_32 ? rules_16_io_n_out_12 : _GEN_282; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_301 = _T_32 ? rules_16_io_n_out_13 : _GEN_283; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_302 = _T_32 ? rules_16_io_n_out_14 : _GEN_284; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_303 = _T_32 ? rules_16_io_n_out_15 : _GEN_285; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_304 = _T_32 ? rules_16_io_n_out_16 : _GEN_286; // @[system.scala 33:21 34:7]
  wire  _GEN_305 = _T_32 ? rules_16_io_x_out : _GEN_287; // @[system.scala 33:21 35:7]
  wire  _T_34 = io_en_a == 7'h11; // @[system.scala 32:27]
  wire [1:0] _GEN_306 = _T_34 ? rules_17_io_n_out_0 : _GEN_288; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_307 = _T_34 ? rules_17_io_n_out_1 : _GEN_289; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_308 = _T_34 ? rules_17_io_n_out_2 : _GEN_290; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_309 = _T_34 ? rules_17_io_n_out_3 : _GEN_291; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_310 = _T_34 ? rules_17_io_n_out_4 : _GEN_292; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_311 = _T_34 ? rules_17_io_n_out_5 : _GEN_293; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_312 = _T_34 ? rules_17_io_n_out_6 : _GEN_294; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_313 = _T_34 ? rules_17_io_n_out_7 : _GEN_295; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_314 = _T_34 ? rules_17_io_n_out_8 : _GEN_296; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_315 = _T_34 ? rules_17_io_n_out_9 : _GEN_297; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_316 = _T_34 ? rules_17_io_n_out_10 : _GEN_298; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_317 = _T_34 ? rules_17_io_n_out_11 : _GEN_299; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_318 = _T_34 ? rules_17_io_n_out_12 : _GEN_300; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_319 = _T_34 ? rules_17_io_n_out_13 : _GEN_301; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_320 = _T_34 ? rules_17_io_n_out_14 : _GEN_302; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_321 = _T_34 ? rules_17_io_n_out_15 : _GEN_303; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_322 = _T_34 ? rules_17_io_n_out_16 : _GEN_304; // @[system.scala 33:21 34:7]
  wire  _GEN_323 = _T_34 ? rules_17_io_x_out : _GEN_305; // @[system.scala 33:21 35:7]
  wire  _T_36 = io_en_a == 7'h12; // @[system.scala 32:27]
  wire [1:0] _GEN_324 = _T_36 ? rules_18_io_n_out_0 : _GEN_306; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_325 = _T_36 ? rules_18_io_n_out_1 : _GEN_307; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_326 = _T_36 ? rules_18_io_n_out_2 : _GEN_308; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_327 = _T_36 ? rules_18_io_n_out_3 : _GEN_309; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_328 = _T_36 ? rules_18_io_n_out_4 : _GEN_310; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_329 = _T_36 ? rules_18_io_n_out_5 : _GEN_311; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_330 = _T_36 ? rules_18_io_n_out_6 : _GEN_312; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_331 = _T_36 ? rules_18_io_n_out_7 : _GEN_313; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_332 = _T_36 ? rules_18_io_n_out_8 : _GEN_314; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_333 = _T_36 ? rules_18_io_n_out_9 : _GEN_315; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_334 = _T_36 ? rules_18_io_n_out_10 : _GEN_316; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_335 = _T_36 ? rules_18_io_n_out_11 : _GEN_317; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_336 = _T_36 ? rules_18_io_n_out_12 : _GEN_318; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_337 = _T_36 ? rules_18_io_n_out_13 : _GEN_319; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_338 = _T_36 ? rules_18_io_n_out_14 : _GEN_320; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_339 = _T_36 ? rules_18_io_n_out_15 : _GEN_321; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_340 = _T_36 ? rules_18_io_n_out_16 : _GEN_322; // @[system.scala 33:21 34:7]
  wire  _GEN_341 = _T_36 ? rules_18_io_x_out : _GEN_323; // @[system.scala 33:21 35:7]
  wire  _T_38 = io_en_a == 7'h13; // @[system.scala 32:27]
  wire [1:0] _GEN_342 = _T_38 ? rules_19_io_n_out_0 : _GEN_324; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_343 = _T_38 ? rules_19_io_n_out_1 : _GEN_325; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_344 = _T_38 ? rules_19_io_n_out_2 : _GEN_326; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_345 = _T_38 ? rules_19_io_n_out_3 : _GEN_327; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_346 = _T_38 ? rules_19_io_n_out_4 : _GEN_328; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_347 = _T_38 ? rules_19_io_n_out_5 : _GEN_329; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_348 = _T_38 ? rules_19_io_n_out_6 : _GEN_330; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_349 = _T_38 ? rules_19_io_n_out_7 : _GEN_331; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_350 = _T_38 ? rules_19_io_n_out_8 : _GEN_332; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_351 = _T_38 ? rules_19_io_n_out_9 : _GEN_333; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_352 = _T_38 ? rules_19_io_n_out_10 : _GEN_334; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_353 = _T_38 ? rules_19_io_n_out_11 : _GEN_335; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_354 = _T_38 ? rules_19_io_n_out_12 : _GEN_336; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_355 = _T_38 ? rules_19_io_n_out_13 : _GEN_337; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_356 = _T_38 ? rules_19_io_n_out_14 : _GEN_338; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_357 = _T_38 ? rules_19_io_n_out_15 : _GEN_339; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_358 = _T_38 ? rules_19_io_n_out_16 : _GEN_340; // @[system.scala 33:21 34:7]
  wire  _GEN_359 = _T_38 ? rules_19_io_x_out : _GEN_341; // @[system.scala 33:21 35:7]
  wire  _T_40 = io_en_a == 7'h14; // @[system.scala 32:27]
  wire [1:0] _GEN_360 = _T_40 ? rules_20_io_n_out_0 : _GEN_342; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_361 = _T_40 ? rules_20_io_n_out_1 : _GEN_343; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_362 = _T_40 ? rules_20_io_n_out_2 : _GEN_344; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_363 = _T_40 ? rules_20_io_n_out_3 : _GEN_345; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_364 = _T_40 ? rules_20_io_n_out_4 : _GEN_346; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_365 = _T_40 ? rules_20_io_n_out_5 : _GEN_347; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_366 = _T_40 ? rules_20_io_n_out_6 : _GEN_348; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_367 = _T_40 ? rules_20_io_n_out_7 : _GEN_349; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_368 = _T_40 ? rules_20_io_n_out_8 : _GEN_350; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_369 = _T_40 ? rules_20_io_n_out_9 : _GEN_351; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_370 = _T_40 ? rules_20_io_n_out_10 : _GEN_352; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_371 = _T_40 ? rules_20_io_n_out_11 : _GEN_353; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_372 = _T_40 ? rules_20_io_n_out_12 : _GEN_354; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_373 = _T_40 ? rules_20_io_n_out_13 : _GEN_355; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_374 = _T_40 ? rules_20_io_n_out_14 : _GEN_356; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_375 = _T_40 ? rules_20_io_n_out_15 : _GEN_357; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_376 = _T_40 ? rules_20_io_n_out_16 : _GEN_358; // @[system.scala 33:21 34:7]
  wire  _GEN_377 = _T_40 ? rules_20_io_x_out : _GEN_359; // @[system.scala 33:21 35:7]
  wire  _T_42 = io_en_a == 7'h15; // @[system.scala 32:27]
  wire [1:0] _GEN_378 = _T_42 ? rules_21_io_n_out_0 : _GEN_360; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_379 = _T_42 ? rules_21_io_n_out_1 : _GEN_361; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_380 = _T_42 ? rules_21_io_n_out_2 : _GEN_362; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_381 = _T_42 ? rules_21_io_n_out_3 : _GEN_363; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_382 = _T_42 ? rules_21_io_n_out_4 : _GEN_364; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_383 = _T_42 ? rules_21_io_n_out_5 : _GEN_365; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_384 = _T_42 ? rules_21_io_n_out_6 : _GEN_366; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_385 = _T_42 ? rules_21_io_n_out_7 : _GEN_367; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_386 = _T_42 ? rules_21_io_n_out_8 : _GEN_368; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_387 = _T_42 ? rules_21_io_n_out_9 : _GEN_369; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_388 = _T_42 ? rules_21_io_n_out_10 : _GEN_370; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_389 = _T_42 ? rules_21_io_n_out_11 : _GEN_371; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_390 = _T_42 ? rules_21_io_n_out_12 : _GEN_372; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_391 = _T_42 ? rules_21_io_n_out_13 : _GEN_373; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_392 = _T_42 ? rules_21_io_n_out_14 : _GEN_374; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_393 = _T_42 ? rules_21_io_n_out_15 : _GEN_375; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_394 = _T_42 ? rules_21_io_n_out_16 : _GEN_376; // @[system.scala 33:21 34:7]
  wire  _GEN_395 = _T_42 ? rules_21_io_x_out : _GEN_377; // @[system.scala 33:21 35:7]
  wire  _T_44 = io_en_a == 7'h16; // @[system.scala 32:27]
  wire [1:0] _GEN_396 = _T_44 ? rules_22_io_n_out_0 : _GEN_378; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_397 = _T_44 ? rules_22_io_n_out_1 : _GEN_379; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_398 = _T_44 ? rules_22_io_n_out_2 : _GEN_380; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_399 = _T_44 ? rules_22_io_n_out_3 : _GEN_381; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_400 = _T_44 ? rules_22_io_n_out_4 : _GEN_382; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_401 = _T_44 ? rules_22_io_n_out_5 : _GEN_383; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_402 = _T_44 ? rules_22_io_n_out_6 : _GEN_384; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_403 = _T_44 ? rules_22_io_n_out_7 : _GEN_385; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_404 = _T_44 ? rules_22_io_n_out_8 : _GEN_386; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_405 = _T_44 ? rules_22_io_n_out_9 : _GEN_387; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_406 = _T_44 ? rules_22_io_n_out_10 : _GEN_388; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_407 = _T_44 ? rules_22_io_n_out_11 : _GEN_389; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_408 = _T_44 ? rules_22_io_n_out_12 : _GEN_390; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_409 = _T_44 ? rules_22_io_n_out_13 : _GEN_391; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_410 = _T_44 ? rules_22_io_n_out_14 : _GEN_392; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_411 = _T_44 ? rules_22_io_n_out_15 : _GEN_393; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_412 = _T_44 ? rules_22_io_n_out_16 : _GEN_394; // @[system.scala 33:21 34:7]
  wire  _GEN_413 = _T_44 ? rules_22_io_x_out : _GEN_395; // @[system.scala 33:21 35:7]
  wire  _T_46 = io_en_a == 7'h17; // @[system.scala 32:27]
  wire [1:0] _GEN_414 = _T_46 ? rules_23_io_n_out_0 : _GEN_396; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_415 = _T_46 ? rules_23_io_n_out_1 : _GEN_397; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_416 = _T_46 ? rules_23_io_n_out_2 : _GEN_398; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_417 = _T_46 ? rules_23_io_n_out_3 : _GEN_399; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_418 = _T_46 ? rules_23_io_n_out_4 : _GEN_400; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_419 = _T_46 ? rules_23_io_n_out_5 : _GEN_401; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_420 = _T_46 ? rules_23_io_n_out_6 : _GEN_402; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_421 = _T_46 ? rules_23_io_n_out_7 : _GEN_403; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_422 = _T_46 ? rules_23_io_n_out_8 : _GEN_404; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_423 = _T_46 ? rules_23_io_n_out_9 : _GEN_405; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_424 = _T_46 ? rules_23_io_n_out_10 : _GEN_406; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_425 = _T_46 ? rules_23_io_n_out_11 : _GEN_407; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_426 = _T_46 ? rules_23_io_n_out_12 : _GEN_408; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_427 = _T_46 ? rules_23_io_n_out_13 : _GEN_409; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_428 = _T_46 ? rules_23_io_n_out_14 : _GEN_410; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_429 = _T_46 ? rules_23_io_n_out_15 : _GEN_411; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_430 = _T_46 ? rules_23_io_n_out_16 : _GEN_412; // @[system.scala 33:21 34:7]
  wire  _GEN_431 = _T_46 ? rules_23_io_x_out : _GEN_413; // @[system.scala 33:21 35:7]
  wire  _T_48 = io_en_a == 7'h18; // @[system.scala 32:27]
  wire [1:0] _GEN_432 = _T_48 ? rules_24_io_n_out_0 : _GEN_414; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_433 = _T_48 ? rules_24_io_n_out_1 : _GEN_415; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_434 = _T_48 ? rules_24_io_n_out_2 : _GEN_416; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_435 = _T_48 ? rules_24_io_n_out_3 : _GEN_417; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_436 = _T_48 ? rules_24_io_n_out_4 : _GEN_418; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_437 = _T_48 ? rules_24_io_n_out_5 : _GEN_419; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_438 = _T_48 ? rules_24_io_n_out_6 : _GEN_420; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_439 = _T_48 ? rules_24_io_n_out_7 : _GEN_421; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_440 = _T_48 ? rules_24_io_n_out_8 : _GEN_422; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_441 = _T_48 ? rules_24_io_n_out_9 : _GEN_423; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_442 = _T_48 ? rules_24_io_n_out_10 : _GEN_424; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_443 = _T_48 ? rules_24_io_n_out_11 : _GEN_425; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_444 = _T_48 ? rules_24_io_n_out_12 : _GEN_426; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_445 = _T_48 ? rules_24_io_n_out_13 : _GEN_427; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_446 = _T_48 ? rules_24_io_n_out_14 : _GEN_428; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_447 = _T_48 ? rules_24_io_n_out_15 : _GEN_429; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_448 = _T_48 ? rules_24_io_n_out_16 : _GEN_430; // @[system.scala 33:21 34:7]
  wire  _GEN_449 = _T_48 ? rules_24_io_x_out : _GEN_431; // @[system.scala 33:21 35:7]
  wire  _T_50 = io_en_a == 7'h19; // @[system.scala 32:27]
  wire [1:0] _GEN_450 = _T_50 ? rules_25_io_n_out_0 : _GEN_432; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_451 = _T_50 ? rules_25_io_n_out_1 : _GEN_433; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_452 = _T_50 ? rules_25_io_n_out_2 : _GEN_434; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_453 = _T_50 ? rules_25_io_n_out_3 : _GEN_435; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_454 = _T_50 ? rules_25_io_n_out_4 : _GEN_436; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_455 = _T_50 ? rules_25_io_n_out_5 : _GEN_437; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_456 = _T_50 ? rules_25_io_n_out_6 : _GEN_438; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_457 = _T_50 ? rules_25_io_n_out_7 : _GEN_439; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_458 = _T_50 ? rules_25_io_n_out_8 : _GEN_440; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_459 = _T_50 ? rules_25_io_n_out_9 : _GEN_441; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_460 = _T_50 ? rules_25_io_n_out_10 : _GEN_442; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_461 = _T_50 ? rules_25_io_n_out_11 : _GEN_443; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_462 = _T_50 ? rules_25_io_n_out_12 : _GEN_444; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_463 = _T_50 ? rules_25_io_n_out_13 : _GEN_445; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_464 = _T_50 ? rules_25_io_n_out_14 : _GEN_446; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_465 = _T_50 ? rules_25_io_n_out_15 : _GEN_447; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_466 = _T_50 ? rules_25_io_n_out_16 : _GEN_448; // @[system.scala 33:21 34:7]
  wire  _GEN_467 = _T_50 ? rules_25_io_x_out : _GEN_449; // @[system.scala 33:21 35:7]
  wire  _T_52 = io_en_a == 7'h1a; // @[system.scala 32:27]
  wire [1:0] _GEN_468 = _T_52 ? rules_26_io_n_out_0 : _GEN_450; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_469 = _T_52 ? rules_26_io_n_out_1 : _GEN_451; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_470 = _T_52 ? rules_26_io_n_out_2 : _GEN_452; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_471 = _T_52 ? rules_26_io_n_out_3 : _GEN_453; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_472 = _T_52 ? rules_26_io_n_out_4 : _GEN_454; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_473 = _T_52 ? rules_26_io_n_out_5 : _GEN_455; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_474 = _T_52 ? rules_26_io_n_out_6 : _GEN_456; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_475 = _T_52 ? rules_26_io_n_out_7 : _GEN_457; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_476 = _T_52 ? rules_26_io_n_out_8 : _GEN_458; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_477 = _T_52 ? rules_26_io_n_out_9 : _GEN_459; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_478 = _T_52 ? rules_26_io_n_out_10 : _GEN_460; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_479 = _T_52 ? rules_26_io_n_out_11 : _GEN_461; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_480 = _T_52 ? rules_26_io_n_out_12 : _GEN_462; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_481 = _T_52 ? rules_26_io_n_out_13 : _GEN_463; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_482 = _T_52 ? rules_26_io_n_out_14 : _GEN_464; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_483 = _T_52 ? rules_26_io_n_out_15 : _GEN_465; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_484 = _T_52 ? rules_26_io_n_out_16 : _GEN_466; // @[system.scala 33:21 34:7]
  wire  _GEN_485 = _T_52 ? rules_26_io_x_out : _GEN_467; // @[system.scala 33:21 35:7]
  wire  _T_54 = io_en_a == 7'h1b; // @[system.scala 32:27]
  wire [1:0] _GEN_486 = _T_54 ? rules_27_io_n_out_0 : _GEN_468; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_487 = _T_54 ? rules_27_io_n_out_1 : _GEN_469; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_488 = _T_54 ? rules_27_io_n_out_2 : _GEN_470; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_489 = _T_54 ? rules_27_io_n_out_3 : _GEN_471; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_490 = _T_54 ? rules_27_io_n_out_4 : _GEN_472; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_491 = _T_54 ? rules_27_io_n_out_5 : _GEN_473; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_492 = _T_54 ? rules_27_io_n_out_6 : _GEN_474; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_493 = _T_54 ? rules_27_io_n_out_7 : _GEN_475; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_494 = _T_54 ? rules_27_io_n_out_8 : _GEN_476; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_495 = _T_54 ? rules_27_io_n_out_9 : _GEN_477; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_496 = _T_54 ? rules_27_io_n_out_10 : _GEN_478; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_497 = _T_54 ? rules_27_io_n_out_11 : _GEN_479; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_498 = _T_54 ? rules_27_io_n_out_12 : _GEN_480; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_499 = _T_54 ? rules_27_io_n_out_13 : _GEN_481; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_500 = _T_54 ? rules_27_io_n_out_14 : _GEN_482; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_501 = _T_54 ? rules_27_io_n_out_15 : _GEN_483; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_502 = _T_54 ? rules_27_io_n_out_16 : _GEN_484; // @[system.scala 33:21 34:7]
  wire  _GEN_503 = _T_54 ? rules_27_io_x_out : _GEN_485; // @[system.scala 33:21 35:7]
  wire  _T_56 = io_en_a == 7'h1c; // @[system.scala 32:27]
  wire [1:0] _GEN_504 = _T_56 ? rules_28_io_n_out_0 : _GEN_486; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_505 = _T_56 ? rules_28_io_n_out_1 : _GEN_487; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_506 = _T_56 ? rules_28_io_n_out_2 : _GEN_488; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_507 = _T_56 ? rules_28_io_n_out_3 : _GEN_489; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_508 = _T_56 ? rules_28_io_n_out_4 : _GEN_490; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_509 = _T_56 ? rules_28_io_n_out_5 : _GEN_491; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_510 = _T_56 ? rules_28_io_n_out_6 : _GEN_492; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_511 = _T_56 ? rules_28_io_n_out_7 : _GEN_493; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_512 = _T_56 ? rules_28_io_n_out_8 : _GEN_494; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_513 = _T_56 ? rules_28_io_n_out_9 : _GEN_495; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_514 = _T_56 ? rules_28_io_n_out_10 : _GEN_496; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_515 = _T_56 ? rules_28_io_n_out_11 : _GEN_497; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_516 = _T_56 ? rules_28_io_n_out_12 : _GEN_498; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_517 = _T_56 ? rules_28_io_n_out_13 : _GEN_499; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_518 = _T_56 ? rules_28_io_n_out_14 : _GEN_500; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_519 = _T_56 ? rules_28_io_n_out_15 : _GEN_501; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_520 = _T_56 ? rules_28_io_n_out_16 : _GEN_502; // @[system.scala 33:21 34:7]
  wire  _GEN_521 = _T_56 ? rules_28_io_x_out : _GEN_503; // @[system.scala 33:21 35:7]
  wire  _T_58 = io_en_a == 7'h1d; // @[system.scala 32:27]
  wire [1:0] _GEN_522 = _T_58 ? rules_29_io_n_out_0 : _GEN_504; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_523 = _T_58 ? rules_29_io_n_out_1 : _GEN_505; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_524 = _T_58 ? rules_29_io_n_out_2 : _GEN_506; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_525 = _T_58 ? rules_29_io_n_out_3 : _GEN_507; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_526 = _T_58 ? rules_29_io_n_out_4 : _GEN_508; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_527 = _T_58 ? rules_29_io_n_out_5 : _GEN_509; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_528 = _T_58 ? rules_29_io_n_out_6 : _GEN_510; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_529 = _T_58 ? rules_29_io_n_out_7 : _GEN_511; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_530 = _T_58 ? rules_29_io_n_out_8 : _GEN_512; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_531 = _T_58 ? rules_29_io_n_out_9 : _GEN_513; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_532 = _T_58 ? rules_29_io_n_out_10 : _GEN_514; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_533 = _T_58 ? rules_29_io_n_out_11 : _GEN_515; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_534 = _T_58 ? rules_29_io_n_out_12 : _GEN_516; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_535 = _T_58 ? rules_29_io_n_out_13 : _GEN_517; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_536 = _T_58 ? rules_29_io_n_out_14 : _GEN_518; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_537 = _T_58 ? rules_29_io_n_out_15 : _GEN_519; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_538 = _T_58 ? rules_29_io_n_out_16 : _GEN_520; // @[system.scala 33:21 34:7]
  wire  _GEN_539 = _T_58 ? rules_29_io_x_out : _GEN_521; // @[system.scala 33:21 35:7]
  wire  _T_60 = io_en_a == 7'h1e; // @[system.scala 32:27]
  wire [1:0] _GEN_540 = _T_60 ? rules_30_io_n_out_0 : _GEN_522; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_541 = _T_60 ? rules_30_io_n_out_1 : _GEN_523; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_542 = _T_60 ? rules_30_io_n_out_2 : _GEN_524; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_543 = _T_60 ? rules_30_io_n_out_3 : _GEN_525; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_544 = _T_60 ? rules_30_io_n_out_4 : _GEN_526; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_545 = _T_60 ? rules_30_io_n_out_5 : _GEN_527; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_546 = _T_60 ? rules_30_io_n_out_6 : _GEN_528; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_547 = _T_60 ? rules_30_io_n_out_7 : _GEN_529; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_548 = _T_60 ? rules_30_io_n_out_8 : _GEN_530; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_549 = _T_60 ? rules_30_io_n_out_9 : _GEN_531; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_550 = _T_60 ? rules_30_io_n_out_10 : _GEN_532; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_551 = _T_60 ? rules_30_io_n_out_11 : _GEN_533; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_552 = _T_60 ? rules_30_io_n_out_12 : _GEN_534; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_553 = _T_60 ? rules_30_io_n_out_13 : _GEN_535; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_554 = _T_60 ? rules_30_io_n_out_14 : _GEN_536; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_555 = _T_60 ? rules_30_io_n_out_15 : _GEN_537; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_556 = _T_60 ? rules_30_io_n_out_16 : _GEN_538; // @[system.scala 33:21 34:7]
  wire  _GEN_557 = _T_60 ? rules_30_io_x_out : _GEN_539; // @[system.scala 33:21 35:7]
  wire  _T_62 = io_en_a == 7'h1f; // @[system.scala 32:27]
  wire [1:0] _GEN_558 = _T_62 ? rules_31_io_n_out_0 : _GEN_540; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_559 = _T_62 ? rules_31_io_n_out_1 : _GEN_541; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_560 = _T_62 ? rules_31_io_n_out_2 : _GEN_542; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_561 = _T_62 ? rules_31_io_n_out_3 : _GEN_543; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_562 = _T_62 ? rules_31_io_n_out_4 : _GEN_544; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_563 = _T_62 ? rules_31_io_n_out_5 : _GEN_545; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_564 = _T_62 ? rules_31_io_n_out_6 : _GEN_546; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_565 = _T_62 ? rules_31_io_n_out_7 : _GEN_547; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_566 = _T_62 ? rules_31_io_n_out_8 : _GEN_548; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_567 = _T_62 ? rules_31_io_n_out_9 : _GEN_549; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_568 = _T_62 ? rules_31_io_n_out_10 : _GEN_550; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_569 = _T_62 ? rules_31_io_n_out_11 : _GEN_551; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_570 = _T_62 ? rules_31_io_n_out_12 : _GEN_552; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_571 = _T_62 ? rules_31_io_n_out_13 : _GEN_553; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_572 = _T_62 ? rules_31_io_n_out_14 : _GEN_554; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_573 = _T_62 ? rules_31_io_n_out_15 : _GEN_555; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_574 = _T_62 ? rules_31_io_n_out_16 : _GEN_556; // @[system.scala 33:21 34:7]
  wire  _GEN_575 = _T_62 ? rules_31_io_x_out : _GEN_557; // @[system.scala 33:21 35:7]
  wire  _T_64 = io_en_a == 7'h20; // @[system.scala 32:27]
  wire [1:0] _GEN_576 = _T_64 ? rules_32_io_n_out_0 : _GEN_558; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_577 = _T_64 ? rules_32_io_n_out_1 : _GEN_559; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_578 = _T_64 ? rules_32_io_n_out_2 : _GEN_560; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_579 = _T_64 ? rules_32_io_n_out_3 : _GEN_561; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_580 = _T_64 ? rules_32_io_n_out_4 : _GEN_562; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_581 = _T_64 ? rules_32_io_n_out_5 : _GEN_563; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_582 = _T_64 ? rules_32_io_n_out_6 : _GEN_564; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_583 = _T_64 ? rules_32_io_n_out_7 : _GEN_565; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_584 = _T_64 ? rules_32_io_n_out_8 : _GEN_566; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_585 = _T_64 ? rules_32_io_n_out_9 : _GEN_567; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_586 = _T_64 ? rules_32_io_n_out_10 : _GEN_568; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_587 = _T_64 ? rules_32_io_n_out_11 : _GEN_569; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_588 = _T_64 ? rules_32_io_n_out_12 : _GEN_570; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_589 = _T_64 ? rules_32_io_n_out_13 : _GEN_571; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_590 = _T_64 ? rules_32_io_n_out_14 : _GEN_572; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_591 = _T_64 ? rules_32_io_n_out_15 : _GEN_573; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_592 = _T_64 ? rules_32_io_n_out_16 : _GEN_574; // @[system.scala 33:21 34:7]
  wire  _GEN_593 = _T_64 ? rules_32_io_x_out : _GEN_575; // @[system.scala 33:21 35:7]
  wire  _T_66 = io_en_a == 7'h21; // @[system.scala 32:27]
  wire [1:0] _GEN_594 = _T_66 ? rules_33_io_n_out_0 : _GEN_576; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_595 = _T_66 ? rules_33_io_n_out_1 : _GEN_577; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_596 = _T_66 ? rules_33_io_n_out_2 : _GEN_578; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_597 = _T_66 ? rules_33_io_n_out_3 : _GEN_579; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_598 = _T_66 ? rules_33_io_n_out_4 : _GEN_580; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_599 = _T_66 ? rules_33_io_n_out_5 : _GEN_581; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_600 = _T_66 ? rules_33_io_n_out_6 : _GEN_582; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_601 = _T_66 ? rules_33_io_n_out_7 : _GEN_583; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_602 = _T_66 ? rules_33_io_n_out_8 : _GEN_584; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_603 = _T_66 ? rules_33_io_n_out_9 : _GEN_585; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_604 = _T_66 ? rules_33_io_n_out_10 : _GEN_586; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_605 = _T_66 ? rules_33_io_n_out_11 : _GEN_587; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_606 = _T_66 ? rules_33_io_n_out_12 : _GEN_588; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_607 = _T_66 ? rules_33_io_n_out_13 : _GEN_589; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_608 = _T_66 ? rules_33_io_n_out_14 : _GEN_590; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_609 = _T_66 ? rules_33_io_n_out_15 : _GEN_591; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_610 = _T_66 ? rules_33_io_n_out_16 : _GEN_592; // @[system.scala 33:21 34:7]
  wire  _GEN_611 = _T_66 ? rules_33_io_x_out : _GEN_593; // @[system.scala 33:21 35:7]
  wire  _T_68 = io_en_a == 7'h22; // @[system.scala 32:27]
  wire [1:0] _GEN_612 = _T_68 ? rules_34_io_n_out_0 : _GEN_594; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_613 = _T_68 ? rules_34_io_n_out_1 : _GEN_595; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_614 = _T_68 ? rules_34_io_n_out_2 : _GEN_596; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_615 = _T_68 ? rules_34_io_n_out_3 : _GEN_597; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_616 = _T_68 ? rules_34_io_n_out_4 : _GEN_598; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_617 = _T_68 ? rules_34_io_n_out_5 : _GEN_599; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_618 = _T_68 ? rules_34_io_n_out_6 : _GEN_600; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_619 = _T_68 ? rules_34_io_n_out_7 : _GEN_601; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_620 = _T_68 ? rules_34_io_n_out_8 : _GEN_602; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_621 = _T_68 ? rules_34_io_n_out_9 : _GEN_603; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_622 = _T_68 ? rules_34_io_n_out_10 : _GEN_604; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_623 = _T_68 ? rules_34_io_n_out_11 : _GEN_605; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_624 = _T_68 ? rules_34_io_n_out_12 : _GEN_606; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_625 = _T_68 ? rules_34_io_n_out_13 : _GEN_607; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_626 = _T_68 ? rules_34_io_n_out_14 : _GEN_608; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_627 = _T_68 ? rules_34_io_n_out_15 : _GEN_609; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_628 = _T_68 ? rules_34_io_n_out_16 : _GEN_610; // @[system.scala 33:21 34:7]
  wire  _GEN_629 = _T_68 ? rules_34_io_x_out : _GEN_611; // @[system.scala 33:21 35:7]
  wire  _T_70 = io_en_a == 7'h23; // @[system.scala 32:27]
  wire [1:0] _GEN_630 = _T_70 ? rules_35_io_n_out_0 : _GEN_612; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_631 = _T_70 ? rules_35_io_n_out_1 : _GEN_613; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_632 = _T_70 ? rules_35_io_n_out_2 : _GEN_614; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_633 = _T_70 ? rules_35_io_n_out_3 : _GEN_615; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_634 = _T_70 ? rules_35_io_n_out_4 : _GEN_616; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_635 = _T_70 ? rules_35_io_n_out_5 : _GEN_617; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_636 = _T_70 ? rules_35_io_n_out_6 : _GEN_618; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_637 = _T_70 ? rules_35_io_n_out_7 : _GEN_619; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_638 = _T_70 ? rules_35_io_n_out_8 : _GEN_620; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_639 = _T_70 ? rules_35_io_n_out_9 : _GEN_621; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_640 = _T_70 ? rules_35_io_n_out_10 : _GEN_622; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_641 = _T_70 ? rules_35_io_n_out_11 : _GEN_623; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_642 = _T_70 ? rules_35_io_n_out_12 : _GEN_624; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_643 = _T_70 ? rules_35_io_n_out_13 : _GEN_625; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_644 = _T_70 ? rules_35_io_n_out_14 : _GEN_626; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_645 = _T_70 ? rules_35_io_n_out_15 : _GEN_627; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_646 = _T_70 ? rules_35_io_n_out_16 : _GEN_628; // @[system.scala 33:21 34:7]
  wire  _GEN_647 = _T_70 ? rules_35_io_x_out : _GEN_629; // @[system.scala 33:21 35:7]
  wire  _T_72 = io_en_a == 7'h24; // @[system.scala 32:27]
  wire [1:0] _GEN_648 = _T_72 ? rules_36_io_n_out_0 : _GEN_630; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_649 = _T_72 ? rules_36_io_n_out_1 : _GEN_631; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_650 = _T_72 ? rules_36_io_n_out_2 : _GEN_632; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_651 = _T_72 ? rules_36_io_n_out_3 : _GEN_633; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_652 = _T_72 ? rules_36_io_n_out_4 : _GEN_634; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_653 = _T_72 ? rules_36_io_n_out_5 : _GEN_635; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_654 = _T_72 ? rules_36_io_n_out_6 : _GEN_636; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_655 = _T_72 ? rules_36_io_n_out_7 : _GEN_637; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_656 = _T_72 ? rules_36_io_n_out_8 : _GEN_638; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_657 = _T_72 ? rules_36_io_n_out_9 : _GEN_639; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_658 = _T_72 ? rules_36_io_n_out_10 : _GEN_640; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_659 = _T_72 ? rules_36_io_n_out_11 : _GEN_641; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_660 = _T_72 ? rules_36_io_n_out_12 : _GEN_642; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_661 = _T_72 ? rules_36_io_n_out_13 : _GEN_643; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_662 = _T_72 ? rules_36_io_n_out_14 : _GEN_644; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_663 = _T_72 ? rules_36_io_n_out_15 : _GEN_645; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_664 = _T_72 ? rules_36_io_n_out_16 : _GEN_646; // @[system.scala 33:21 34:7]
  wire  _GEN_665 = _T_72 ? rules_36_io_x_out : _GEN_647; // @[system.scala 33:21 35:7]
  wire  _T_74 = io_en_a == 7'h25; // @[system.scala 32:27]
  wire [1:0] _GEN_666 = _T_74 ? rules_37_io_n_out_0 : _GEN_648; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_667 = _T_74 ? rules_37_io_n_out_1 : _GEN_649; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_668 = _T_74 ? rules_37_io_n_out_2 : _GEN_650; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_669 = _T_74 ? rules_37_io_n_out_3 : _GEN_651; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_670 = _T_74 ? rules_37_io_n_out_4 : _GEN_652; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_671 = _T_74 ? rules_37_io_n_out_5 : _GEN_653; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_672 = _T_74 ? rules_37_io_n_out_6 : _GEN_654; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_673 = _T_74 ? rules_37_io_n_out_7 : _GEN_655; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_674 = _T_74 ? rules_37_io_n_out_8 : _GEN_656; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_675 = _T_74 ? rules_37_io_n_out_9 : _GEN_657; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_676 = _T_74 ? rules_37_io_n_out_10 : _GEN_658; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_677 = _T_74 ? rules_37_io_n_out_11 : _GEN_659; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_678 = _T_74 ? rules_37_io_n_out_12 : _GEN_660; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_679 = _T_74 ? rules_37_io_n_out_13 : _GEN_661; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_680 = _T_74 ? rules_37_io_n_out_14 : _GEN_662; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_681 = _T_74 ? rules_37_io_n_out_15 : _GEN_663; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_682 = _T_74 ? rules_37_io_n_out_16 : _GEN_664; // @[system.scala 33:21 34:7]
  wire  _GEN_683 = _T_74 ? rules_37_io_x_out : _GEN_665; // @[system.scala 33:21 35:7]
  wire  _T_76 = io_en_a == 7'h26; // @[system.scala 32:27]
  wire [1:0] _GEN_684 = _T_76 ? rules_38_io_n_out_0 : _GEN_666; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_685 = _T_76 ? rules_38_io_n_out_1 : _GEN_667; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_686 = _T_76 ? rules_38_io_n_out_2 : _GEN_668; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_687 = _T_76 ? rules_38_io_n_out_3 : _GEN_669; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_688 = _T_76 ? rules_38_io_n_out_4 : _GEN_670; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_689 = _T_76 ? rules_38_io_n_out_5 : _GEN_671; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_690 = _T_76 ? rules_38_io_n_out_6 : _GEN_672; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_691 = _T_76 ? rules_38_io_n_out_7 : _GEN_673; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_692 = _T_76 ? rules_38_io_n_out_8 : _GEN_674; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_693 = _T_76 ? rules_38_io_n_out_9 : _GEN_675; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_694 = _T_76 ? rules_38_io_n_out_10 : _GEN_676; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_695 = _T_76 ? rules_38_io_n_out_11 : _GEN_677; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_696 = _T_76 ? rules_38_io_n_out_12 : _GEN_678; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_697 = _T_76 ? rules_38_io_n_out_13 : _GEN_679; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_698 = _T_76 ? rules_38_io_n_out_14 : _GEN_680; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_699 = _T_76 ? rules_38_io_n_out_15 : _GEN_681; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_700 = _T_76 ? rules_38_io_n_out_16 : _GEN_682; // @[system.scala 33:21 34:7]
  wire  _GEN_701 = _T_76 ? rules_38_io_x_out : _GEN_683; // @[system.scala 33:21 35:7]
  wire  _T_78 = io_en_a == 7'h27; // @[system.scala 32:27]
  wire [1:0] _GEN_702 = _T_78 ? rules_39_io_n_out_0 : _GEN_684; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_703 = _T_78 ? rules_39_io_n_out_1 : _GEN_685; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_704 = _T_78 ? rules_39_io_n_out_2 : _GEN_686; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_705 = _T_78 ? rules_39_io_n_out_3 : _GEN_687; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_706 = _T_78 ? rules_39_io_n_out_4 : _GEN_688; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_707 = _T_78 ? rules_39_io_n_out_5 : _GEN_689; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_708 = _T_78 ? rules_39_io_n_out_6 : _GEN_690; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_709 = _T_78 ? rules_39_io_n_out_7 : _GEN_691; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_710 = _T_78 ? rules_39_io_n_out_8 : _GEN_692; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_711 = _T_78 ? rules_39_io_n_out_9 : _GEN_693; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_712 = _T_78 ? rules_39_io_n_out_10 : _GEN_694; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_713 = _T_78 ? rules_39_io_n_out_11 : _GEN_695; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_714 = _T_78 ? rules_39_io_n_out_12 : _GEN_696; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_715 = _T_78 ? rules_39_io_n_out_13 : _GEN_697; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_716 = _T_78 ? rules_39_io_n_out_14 : _GEN_698; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_717 = _T_78 ? rules_39_io_n_out_15 : _GEN_699; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_718 = _T_78 ? rules_39_io_n_out_16 : _GEN_700; // @[system.scala 33:21 34:7]
  wire  _GEN_719 = _T_78 ? rules_39_io_x_out : _GEN_701; // @[system.scala 33:21 35:7]
  wire  _T_80 = io_en_a == 7'h28; // @[system.scala 32:27]
  wire [1:0] _GEN_720 = _T_80 ? rules_40_io_n_out_0 : _GEN_702; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_721 = _T_80 ? rules_40_io_n_out_1 : _GEN_703; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_722 = _T_80 ? rules_40_io_n_out_2 : _GEN_704; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_723 = _T_80 ? rules_40_io_n_out_3 : _GEN_705; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_724 = _T_80 ? rules_40_io_n_out_4 : _GEN_706; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_725 = _T_80 ? rules_40_io_n_out_5 : _GEN_707; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_726 = _T_80 ? rules_40_io_n_out_6 : _GEN_708; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_727 = _T_80 ? rules_40_io_n_out_7 : _GEN_709; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_728 = _T_80 ? rules_40_io_n_out_8 : _GEN_710; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_729 = _T_80 ? rules_40_io_n_out_9 : _GEN_711; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_730 = _T_80 ? rules_40_io_n_out_10 : _GEN_712; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_731 = _T_80 ? rules_40_io_n_out_11 : _GEN_713; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_732 = _T_80 ? rules_40_io_n_out_12 : _GEN_714; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_733 = _T_80 ? rules_40_io_n_out_13 : _GEN_715; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_734 = _T_80 ? rules_40_io_n_out_14 : _GEN_716; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_735 = _T_80 ? rules_40_io_n_out_15 : _GEN_717; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_736 = _T_80 ? rules_40_io_n_out_16 : _GEN_718; // @[system.scala 33:21 34:7]
  wire  _GEN_737 = _T_80 ? rules_40_io_x_out : _GEN_719; // @[system.scala 33:21 35:7]
  wire  _T_82 = io_en_a == 7'h29; // @[system.scala 32:27]
  wire [1:0] _GEN_738 = _T_82 ? rules_41_io_n_out_0 : _GEN_720; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_739 = _T_82 ? rules_41_io_n_out_1 : _GEN_721; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_740 = _T_82 ? rules_41_io_n_out_2 : _GEN_722; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_741 = _T_82 ? rules_41_io_n_out_3 : _GEN_723; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_742 = _T_82 ? rules_41_io_n_out_4 : _GEN_724; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_743 = _T_82 ? rules_41_io_n_out_5 : _GEN_725; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_744 = _T_82 ? rules_41_io_n_out_6 : _GEN_726; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_745 = _T_82 ? rules_41_io_n_out_7 : _GEN_727; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_746 = _T_82 ? rules_41_io_n_out_8 : _GEN_728; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_747 = _T_82 ? rules_41_io_n_out_9 : _GEN_729; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_748 = _T_82 ? rules_41_io_n_out_10 : _GEN_730; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_749 = _T_82 ? rules_41_io_n_out_11 : _GEN_731; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_750 = _T_82 ? rules_41_io_n_out_12 : _GEN_732; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_751 = _T_82 ? rules_41_io_n_out_13 : _GEN_733; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_752 = _T_82 ? rules_41_io_n_out_14 : _GEN_734; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_753 = _T_82 ? rules_41_io_n_out_15 : _GEN_735; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_754 = _T_82 ? rules_41_io_n_out_16 : _GEN_736; // @[system.scala 33:21 34:7]
  wire  _GEN_755 = _T_82 ? rules_41_io_x_out : _GEN_737; // @[system.scala 33:21 35:7]
  wire  _T_84 = io_en_a == 7'h2a; // @[system.scala 32:27]
  wire [1:0] _GEN_756 = _T_84 ? rules_42_io_n_out_0 : _GEN_738; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_757 = _T_84 ? rules_42_io_n_out_1 : _GEN_739; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_758 = _T_84 ? rules_42_io_n_out_2 : _GEN_740; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_759 = _T_84 ? rules_42_io_n_out_3 : _GEN_741; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_760 = _T_84 ? rules_42_io_n_out_4 : _GEN_742; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_761 = _T_84 ? rules_42_io_n_out_5 : _GEN_743; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_762 = _T_84 ? rules_42_io_n_out_6 : _GEN_744; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_763 = _T_84 ? rules_42_io_n_out_7 : _GEN_745; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_764 = _T_84 ? rules_42_io_n_out_8 : _GEN_746; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_765 = _T_84 ? rules_42_io_n_out_9 : _GEN_747; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_766 = _T_84 ? rules_42_io_n_out_10 : _GEN_748; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_767 = _T_84 ? rules_42_io_n_out_11 : _GEN_749; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_768 = _T_84 ? rules_42_io_n_out_12 : _GEN_750; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_769 = _T_84 ? rules_42_io_n_out_13 : _GEN_751; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_770 = _T_84 ? rules_42_io_n_out_14 : _GEN_752; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_771 = _T_84 ? rules_42_io_n_out_15 : _GEN_753; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_772 = _T_84 ? rules_42_io_n_out_16 : _GEN_754; // @[system.scala 33:21 34:7]
  wire  _GEN_773 = _T_84 ? rules_42_io_x_out : _GEN_755; // @[system.scala 33:21 35:7]
  wire  _T_86 = io_en_a == 7'h2b; // @[system.scala 32:27]
  wire [1:0] _GEN_774 = _T_86 ? rules_43_io_n_out_0 : _GEN_756; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_775 = _T_86 ? rules_43_io_n_out_1 : _GEN_757; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_776 = _T_86 ? rules_43_io_n_out_2 : _GEN_758; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_777 = _T_86 ? rules_43_io_n_out_3 : _GEN_759; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_778 = _T_86 ? rules_43_io_n_out_4 : _GEN_760; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_779 = _T_86 ? rules_43_io_n_out_5 : _GEN_761; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_780 = _T_86 ? rules_43_io_n_out_6 : _GEN_762; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_781 = _T_86 ? rules_43_io_n_out_7 : _GEN_763; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_782 = _T_86 ? rules_43_io_n_out_8 : _GEN_764; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_783 = _T_86 ? rules_43_io_n_out_9 : _GEN_765; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_784 = _T_86 ? rules_43_io_n_out_10 : _GEN_766; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_785 = _T_86 ? rules_43_io_n_out_11 : _GEN_767; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_786 = _T_86 ? rules_43_io_n_out_12 : _GEN_768; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_787 = _T_86 ? rules_43_io_n_out_13 : _GEN_769; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_788 = _T_86 ? rules_43_io_n_out_14 : _GEN_770; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_789 = _T_86 ? rules_43_io_n_out_15 : _GEN_771; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_790 = _T_86 ? rules_43_io_n_out_16 : _GEN_772; // @[system.scala 33:21 34:7]
  wire  _GEN_791 = _T_86 ? rules_43_io_x_out : _GEN_773; // @[system.scala 33:21 35:7]
  wire  _T_88 = io_en_a == 7'h2c; // @[system.scala 32:27]
  wire [1:0] _GEN_792 = _T_88 ? rules_44_io_n_out_0 : _GEN_774; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_793 = _T_88 ? rules_44_io_n_out_1 : _GEN_775; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_794 = _T_88 ? rules_44_io_n_out_2 : _GEN_776; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_795 = _T_88 ? rules_44_io_n_out_3 : _GEN_777; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_796 = _T_88 ? rules_44_io_n_out_4 : _GEN_778; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_797 = _T_88 ? rules_44_io_n_out_5 : _GEN_779; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_798 = _T_88 ? rules_44_io_n_out_6 : _GEN_780; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_799 = _T_88 ? rules_44_io_n_out_7 : _GEN_781; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_800 = _T_88 ? rules_44_io_n_out_8 : _GEN_782; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_801 = _T_88 ? rules_44_io_n_out_9 : _GEN_783; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_802 = _T_88 ? rules_44_io_n_out_10 : _GEN_784; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_803 = _T_88 ? rules_44_io_n_out_11 : _GEN_785; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_804 = _T_88 ? rules_44_io_n_out_12 : _GEN_786; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_805 = _T_88 ? rules_44_io_n_out_13 : _GEN_787; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_806 = _T_88 ? rules_44_io_n_out_14 : _GEN_788; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_807 = _T_88 ? rules_44_io_n_out_15 : _GEN_789; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_808 = _T_88 ? rules_44_io_n_out_16 : _GEN_790; // @[system.scala 33:21 34:7]
  wire  _GEN_809 = _T_88 ? rules_44_io_x_out : _GEN_791; // @[system.scala 33:21 35:7]
  wire  _T_90 = io_en_a == 7'h2d; // @[system.scala 32:27]
  wire [1:0] _GEN_810 = _T_90 ? rules_45_io_n_out_0 : _GEN_792; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_811 = _T_90 ? rules_45_io_n_out_1 : _GEN_793; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_812 = _T_90 ? rules_45_io_n_out_2 : _GEN_794; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_813 = _T_90 ? rules_45_io_n_out_3 : _GEN_795; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_814 = _T_90 ? rules_45_io_n_out_4 : _GEN_796; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_815 = _T_90 ? rules_45_io_n_out_5 : _GEN_797; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_816 = _T_90 ? rules_45_io_n_out_6 : _GEN_798; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_817 = _T_90 ? rules_45_io_n_out_7 : _GEN_799; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_818 = _T_90 ? rules_45_io_n_out_8 : _GEN_800; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_819 = _T_90 ? rules_45_io_n_out_9 : _GEN_801; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_820 = _T_90 ? rules_45_io_n_out_10 : _GEN_802; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_821 = _T_90 ? rules_45_io_n_out_11 : _GEN_803; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_822 = _T_90 ? rules_45_io_n_out_12 : _GEN_804; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_823 = _T_90 ? rules_45_io_n_out_13 : _GEN_805; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_824 = _T_90 ? rules_45_io_n_out_14 : _GEN_806; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_825 = _T_90 ? rules_45_io_n_out_15 : _GEN_807; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_826 = _T_90 ? rules_45_io_n_out_16 : _GEN_808; // @[system.scala 33:21 34:7]
  wire  _GEN_827 = _T_90 ? rules_45_io_x_out : _GEN_809; // @[system.scala 33:21 35:7]
  wire  _T_92 = io_en_a == 7'h2e; // @[system.scala 32:27]
  wire [1:0] _GEN_828 = _T_92 ? rules_46_io_n_out_0 : _GEN_810; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_829 = _T_92 ? rules_46_io_n_out_1 : _GEN_811; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_830 = _T_92 ? rules_46_io_n_out_2 : _GEN_812; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_831 = _T_92 ? rules_46_io_n_out_3 : _GEN_813; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_832 = _T_92 ? rules_46_io_n_out_4 : _GEN_814; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_833 = _T_92 ? rules_46_io_n_out_5 : _GEN_815; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_834 = _T_92 ? rules_46_io_n_out_6 : _GEN_816; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_835 = _T_92 ? rules_46_io_n_out_7 : _GEN_817; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_836 = _T_92 ? rules_46_io_n_out_8 : _GEN_818; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_837 = _T_92 ? rules_46_io_n_out_9 : _GEN_819; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_838 = _T_92 ? rules_46_io_n_out_10 : _GEN_820; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_839 = _T_92 ? rules_46_io_n_out_11 : _GEN_821; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_840 = _T_92 ? rules_46_io_n_out_12 : _GEN_822; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_841 = _T_92 ? rules_46_io_n_out_13 : _GEN_823; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_842 = _T_92 ? rules_46_io_n_out_14 : _GEN_824; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_843 = _T_92 ? rules_46_io_n_out_15 : _GEN_825; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_844 = _T_92 ? rules_46_io_n_out_16 : _GEN_826; // @[system.scala 33:21 34:7]
  wire  _GEN_845 = _T_92 ? rules_46_io_x_out : _GEN_827; // @[system.scala 33:21 35:7]
  wire  _T_94 = io_en_a == 7'h2f; // @[system.scala 32:27]
  wire [1:0] _GEN_846 = _T_94 ? rules_47_io_n_out_0 : _GEN_828; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_847 = _T_94 ? rules_47_io_n_out_1 : _GEN_829; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_848 = _T_94 ? rules_47_io_n_out_2 : _GEN_830; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_849 = _T_94 ? rules_47_io_n_out_3 : _GEN_831; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_850 = _T_94 ? rules_47_io_n_out_4 : _GEN_832; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_851 = _T_94 ? rules_47_io_n_out_5 : _GEN_833; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_852 = _T_94 ? rules_47_io_n_out_6 : _GEN_834; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_853 = _T_94 ? rules_47_io_n_out_7 : _GEN_835; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_854 = _T_94 ? rules_47_io_n_out_8 : _GEN_836; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_855 = _T_94 ? rules_47_io_n_out_9 : _GEN_837; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_856 = _T_94 ? rules_47_io_n_out_10 : _GEN_838; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_857 = _T_94 ? rules_47_io_n_out_11 : _GEN_839; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_858 = _T_94 ? rules_47_io_n_out_12 : _GEN_840; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_859 = _T_94 ? rules_47_io_n_out_13 : _GEN_841; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_860 = _T_94 ? rules_47_io_n_out_14 : _GEN_842; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_861 = _T_94 ? rules_47_io_n_out_15 : _GEN_843; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_862 = _T_94 ? rules_47_io_n_out_16 : _GEN_844; // @[system.scala 33:21 34:7]
  wire  _GEN_863 = _T_94 ? rules_47_io_x_out : _GEN_845; // @[system.scala 33:21 35:7]
  wire  _T_96 = io_en_a == 7'h30; // @[system.scala 32:27]
  wire [1:0] _GEN_864 = _T_96 ? rules_48_io_n_out_0 : _GEN_846; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_865 = _T_96 ? rules_48_io_n_out_1 : _GEN_847; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_866 = _T_96 ? rules_48_io_n_out_2 : _GEN_848; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_867 = _T_96 ? rules_48_io_n_out_3 : _GEN_849; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_868 = _T_96 ? rules_48_io_n_out_4 : _GEN_850; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_869 = _T_96 ? rules_48_io_n_out_5 : _GEN_851; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_870 = _T_96 ? rules_48_io_n_out_6 : _GEN_852; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_871 = _T_96 ? rules_48_io_n_out_7 : _GEN_853; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_872 = _T_96 ? rules_48_io_n_out_8 : _GEN_854; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_873 = _T_96 ? rules_48_io_n_out_9 : _GEN_855; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_874 = _T_96 ? rules_48_io_n_out_10 : _GEN_856; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_875 = _T_96 ? rules_48_io_n_out_11 : _GEN_857; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_876 = _T_96 ? rules_48_io_n_out_12 : _GEN_858; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_877 = _T_96 ? rules_48_io_n_out_13 : _GEN_859; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_878 = _T_96 ? rules_48_io_n_out_14 : _GEN_860; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_879 = _T_96 ? rules_48_io_n_out_15 : _GEN_861; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_880 = _T_96 ? rules_48_io_n_out_16 : _GEN_862; // @[system.scala 33:21 34:7]
  wire  _GEN_881 = _T_96 ? rules_48_io_x_out : _GEN_863; // @[system.scala 33:21 35:7]
  wire  _T_98 = io_en_a == 7'h31; // @[system.scala 32:27]
  wire [1:0] _GEN_882 = _T_98 ? rules_49_io_n_out_0 : _GEN_864; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_883 = _T_98 ? rules_49_io_n_out_1 : _GEN_865; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_884 = _T_98 ? rules_49_io_n_out_2 : _GEN_866; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_885 = _T_98 ? rules_49_io_n_out_3 : _GEN_867; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_886 = _T_98 ? rules_49_io_n_out_4 : _GEN_868; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_887 = _T_98 ? rules_49_io_n_out_5 : _GEN_869; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_888 = _T_98 ? rules_49_io_n_out_6 : _GEN_870; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_889 = _T_98 ? rules_49_io_n_out_7 : _GEN_871; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_890 = _T_98 ? rules_49_io_n_out_8 : _GEN_872; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_891 = _T_98 ? rules_49_io_n_out_9 : _GEN_873; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_892 = _T_98 ? rules_49_io_n_out_10 : _GEN_874; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_893 = _T_98 ? rules_49_io_n_out_11 : _GEN_875; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_894 = _T_98 ? rules_49_io_n_out_12 : _GEN_876; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_895 = _T_98 ? rules_49_io_n_out_13 : _GEN_877; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_896 = _T_98 ? rules_49_io_n_out_14 : _GEN_878; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_897 = _T_98 ? rules_49_io_n_out_15 : _GEN_879; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_898 = _T_98 ? rules_49_io_n_out_16 : _GEN_880; // @[system.scala 33:21 34:7]
  wire  _GEN_899 = _T_98 ? rules_49_io_x_out : _GEN_881; // @[system.scala 33:21 35:7]
  wire  _T_100 = io_en_a == 7'h32; // @[system.scala 32:27]
  wire [1:0] _GEN_900 = _T_100 ? rules_50_io_n_out_0 : _GEN_882; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_901 = _T_100 ? rules_50_io_n_out_1 : _GEN_883; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_902 = _T_100 ? rules_50_io_n_out_2 : _GEN_884; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_903 = _T_100 ? rules_50_io_n_out_3 : _GEN_885; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_904 = _T_100 ? rules_50_io_n_out_4 : _GEN_886; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_905 = _T_100 ? rules_50_io_n_out_5 : _GEN_887; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_906 = _T_100 ? rules_50_io_n_out_6 : _GEN_888; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_907 = _T_100 ? rules_50_io_n_out_7 : _GEN_889; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_908 = _T_100 ? rules_50_io_n_out_8 : _GEN_890; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_909 = _T_100 ? rules_50_io_n_out_9 : _GEN_891; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_910 = _T_100 ? rules_50_io_n_out_10 : _GEN_892; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_911 = _T_100 ? rules_50_io_n_out_11 : _GEN_893; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_912 = _T_100 ? rules_50_io_n_out_12 : _GEN_894; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_913 = _T_100 ? rules_50_io_n_out_13 : _GEN_895; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_914 = _T_100 ? rules_50_io_n_out_14 : _GEN_896; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_915 = _T_100 ? rules_50_io_n_out_15 : _GEN_897; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_916 = _T_100 ? rules_50_io_n_out_16 : _GEN_898; // @[system.scala 33:21 34:7]
  wire  _GEN_917 = _T_100 ? rules_50_io_x_out : _GEN_899; // @[system.scala 33:21 35:7]
  wire  _T_102 = io_en_a == 7'h33; // @[system.scala 32:27]
  wire [1:0] _GEN_918 = _T_102 ? rules_51_io_n_out_0 : _GEN_900; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_919 = _T_102 ? rules_51_io_n_out_1 : _GEN_901; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_920 = _T_102 ? rules_51_io_n_out_2 : _GEN_902; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_921 = _T_102 ? rules_51_io_n_out_3 : _GEN_903; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_922 = _T_102 ? rules_51_io_n_out_4 : _GEN_904; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_923 = _T_102 ? rules_51_io_n_out_5 : _GEN_905; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_924 = _T_102 ? rules_51_io_n_out_6 : _GEN_906; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_925 = _T_102 ? rules_51_io_n_out_7 : _GEN_907; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_926 = _T_102 ? rules_51_io_n_out_8 : _GEN_908; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_927 = _T_102 ? rules_51_io_n_out_9 : _GEN_909; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_928 = _T_102 ? rules_51_io_n_out_10 : _GEN_910; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_929 = _T_102 ? rules_51_io_n_out_11 : _GEN_911; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_930 = _T_102 ? rules_51_io_n_out_12 : _GEN_912; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_931 = _T_102 ? rules_51_io_n_out_13 : _GEN_913; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_932 = _T_102 ? rules_51_io_n_out_14 : _GEN_914; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_933 = _T_102 ? rules_51_io_n_out_15 : _GEN_915; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_934 = _T_102 ? rules_51_io_n_out_16 : _GEN_916; // @[system.scala 33:21 34:7]
  wire  _GEN_935 = _T_102 ? rules_51_io_x_out : _GEN_917; // @[system.scala 33:21 35:7]
  wire  _T_104 = io_en_a == 7'h34; // @[system.scala 32:27]
  wire [1:0] _GEN_936 = _T_104 ? rules_52_io_n_out_0 : _GEN_918; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_937 = _T_104 ? rules_52_io_n_out_1 : _GEN_919; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_938 = _T_104 ? rules_52_io_n_out_2 : _GEN_920; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_939 = _T_104 ? rules_52_io_n_out_3 : _GEN_921; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_940 = _T_104 ? rules_52_io_n_out_4 : _GEN_922; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_941 = _T_104 ? rules_52_io_n_out_5 : _GEN_923; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_942 = _T_104 ? rules_52_io_n_out_6 : _GEN_924; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_943 = _T_104 ? rules_52_io_n_out_7 : _GEN_925; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_944 = _T_104 ? rules_52_io_n_out_8 : _GEN_926; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_945 = _T_104 ? rules_52_io_n_out_9 : _GEN_927; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_946 = _T_104 ? rules_52_io_n_out_10 : _GEN_928; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_947 = _T_104 ? rules_52_io_n_out_11 : _GEN_929; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_948 = _T_104 ? rules_52_io_n_out_12 : _GEN_930; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_949 = _T_104 ? rules_52_io_n_out_13 : _GEN_931; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_950 = _T_104 ? rules_52_io_n_out_14 : _GEN_932; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_951 = _T_104 ? rules_52_io_n_out_15 : _GEN_933; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_952 = _T_104 ? rules_52_io_n_out_16 : _GEN_934; // @[system.scala 33:21 34:7]
  wire  _GEN_953 = _T_104 ? rules_52_io_x_out : _GEN_935; // @[system.scala 33:21 35:7]
  wire  _T_106 = io_en_a == 7'h35; // @[system.scala 32:27]
  wire [1:0] _GEN_954 = _T_106 ? rules_53_io_n_out_0 : _GEN_936; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_955 = _T_106 ? rules_53_io_n_out_1 : _GEN_937; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_956 = _T_106 ? rules_53_io_n_out_2 : _GEN_938; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_957 = _T_106 ? rules_53_io_n_out_3 : _GEN_939; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_958 = _T_106 ? rules_53_io_n_out_4 : _GEN_940; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_959 = _T_106 ? rules_53_io_n_out_5 : _GEN_941; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_960 = _T_106 ? rules_53_io_n_out_6 : _GEN_942; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_961 = _T_106 ? rules_53_io_n_out_7 : _GEN_943; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_962 = _T_106 ? rules_53_io_n_out_8 : _GEN_944; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_963 = _T_106 ? rules_53_io_n_out_9 : _GEN_945; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_964 = _T_106 ? rules_53_io_n_out_10 : _GEN_946; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_965 = _T_106 ? rules_53_io_n_out_11 : _GEN_947; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_966 = _T_106 ? rules_53_io_n_out_12 : _GEN_948; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_967 = _T_106 ? rules_53_io_n_out_13 : _GEN_949; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_968 = _T_106 ? rules_53_io_n_out_14 : _GEN_950; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_969 = _T_106 ? rules_53_io_n_out_15 : _GEN_951; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_970 = _T_106 ? rules_53_io_n_out_16 : _GEN_952; // @[system.scala 33:21 34:7]
  wire  _GEN_971 = _T_106 ? rules_53_io_x_out : _GEN_953; // @[system.scala 33:21 35:7]
  wire  _T_108 = io_en_a == 7'h36; // @[system.scala 32:27]
  wire [1:0] _GEN_972 = _T_108 ? rules_54_io_n_out_0 : _GEN_954; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_973 = _T_108 ? rules_54_io_n_out_1 : _GEN_955; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_974 = _T_108 ? rules_54_io_n_out_2 : _GEN_956; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_975 = _T_108 ? rules_54_io_n_out_3 : _GEN_957; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_976 = _T_108 ? rules_54_io_n_out_4 : _GEN_958; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_977 = _T_108 ? rules_54_io_n_out_5 : _GEN_959; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_978 = _T_108 ? rules_54_io_n_out_6 : _GEN_960; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_979 = _T_108 ? rules_54_io_n_out_7 : _GEN_961; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_980 = _T_108 ? rules_54_io_n_out_8 : _GEN_962; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_981 = _T_108 ? rules_54_io_n_out_9 : _GEN_963; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_982 = _T_108 ? rules_54_io_n_out_10 : _GEN_964; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_983 = _T_108 ? rules_54_io_n_out_11 : _GEN_965; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_984 = _T_108 ? rules_54_io_n_out_12 : _GEN_966; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_985 = _T_108 ? rules_54_io_n_out_13 : _GEN_967; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_986 = _T_108 ? rules_54_io_n_out_14 : _GEN_968; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_987 = _T_108 ? rules_54_io_n_out_15 : _GEN_969; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_988 = _T_108 ? rules_54_io_n_out_16 : _GEN_970; // @[system.scala 33:21 34:7]
  wire  _GEN_989 = _T_108 ? rules_54_io_x_out : _GEN_971; // @[system.scala 33:21 35:7]
  wire  _T_110 = io_en_a == 7'h37; // @[system.scala 32:27]
  wire [1:0] _GEN_990 = _T_110 ? rules_55_io_n_out_0 : _GEN_972; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_991 = _T_110 ? rules_55_io_n_out_1 : _GEN_973; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_992 = _T_110 ? rules_55_io_n_out_2 : _GEN_974; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_993 = _T_110 ? rules_55_io_n_out_3 : _GEN_975; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_994 = _T_110 ? rules_55_io_n_out_4 : _GEN_976; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_995 = _T_110 ? rules_55_io_n_out_5 : _GEN_977; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_996 = _T_110 ? rules_55_io_n_out_6 : _GEN_978; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_997 = _T_110 ? rules_55_io_n_out_7 : _GEN_979; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_998 = _T_110 ? rules_55_io_n_out_8 : _GEN_980; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_999 = _T_110 ? rules_55_io_n_out_9 : _GEN_981; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1000 = _T_110 ? rules_55_io_n_out_10 : _GEN_982; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1001 = _T_110 ? rules_55_io_n_out_11 : _GEN_983; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1002 = _T_110 ? rules_55_io_n_out_12 : _GEN_984; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1003 = _T_110 ? rules_55_io_n_out_13 : _GEN_985; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1004 = _T_110 ? rules_55_io_n_out_14 : _GEN_986; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1005 = _T_110 ? rules_55_io_n_out_15 : _GEN_987; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1006 = _T_110 ? rules_55_io_n_out_16 : _GEN_988; // @[system.scala 33:21 34:7]
  wire  _GEN_1007 = _T_110 ? rules_55_io_x_out : _GEN_989; // @[system.scala 33:21 35:7]
  wire  _T_112 = io_en_a == 7'h38; // @[system.scala 32:27]
  wire [1:0] _GEN_1008 = _T_112 ? rules_56_io_n_out_0 : _GEN_990; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1009 = _T_112 ? rules_56_io_n_out_1 : _GEN_991; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1010 = _T_112 ? rules_56_io_n_out_2 : _GEN_992; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1011 = _T_112 ? rules_56_io_n_out_3 : _GEN_993; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1012 = _T_112 ? rules_56_io_n_out_4 : _GEN_994; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1013 = _T_112 ? rules_56_io_n_out_5 : _GEN_995; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1014 = _T_112 ? rules_56_io_n_out_6 : _GEN_996; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1015 = _T_112 ? rules_56_io_n_out_7 : _GEN_997; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1016 = _T_112 ? rules_56_io_n_out_8 : _GEN_998; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1017 = _T_112 ? rules_56_io_n_out_9 : _GEN_999; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1018 = _T_112 ? rules_56_io_n_out_10 : _GEN_1000; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1019 = _T_112 ? rules_56_io_n_out_11 : _GEN_1001; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1020 = _T_112 ? rules_56_io_n_out_12 : _GEN_1002; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1021 = _T_112 ? rules_56_io_n_out_13 : _GEN_1003; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1022 = _T_112 ? rules_56_io_n_out_14 : _GEN_1004; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1023 = _T_112 ? rules_56_io_n_out_15 : _GEN_1005; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1024 = _T_112 ? rules_56_io_n_out_16 : _GEN_1006; // @[system.scala 33:21 34:7]
  wire  _GEN_1025 = _T_112 ? rules_56_io_x_out : _GEN_1007; // @[system.scala 33:21 35:7]
  wire  _T_114 = io_en_a == 7'h39; // @[system.scala 32:27]
  wire [1:0] _GEN_1026 = _T_114 ? rules_57_io_n_out_0 : _GEN_1008; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1027 = _T_114 ? rules_57_io_n_out_1 : _GEN_1009; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1028 = _T_114 ? rules_57_io_n_out_2 : _GEN_1010; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1029 = _T_114 ? rules_57_io_n_out_3 : _GEN_1011; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1030 = _T_114 ? rules_57_io_n_out_4 : _GEN_1012; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1031 = _T_114 ? rules_57_io_n_out_5 : _GEN_1013; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1032 = _T_114 ? rules_57_io_n_out_6 : _GEN_1014; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1033 = _T_114 ? rules_57_io_n_out_7 : _GEN_1015; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1034 = _T_114 ? rules_57_io_n_out_8 : _GEN_1016; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1035 = _T_114 ? rules_57_io_n_out_9 : _GEN_1017; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1036 = _T_114 ? rules_57_io_n_out_10 : _GEN_1018; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1037 = _T_114 ? rules_57_io_n_out_11 : _GEN_1019; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1038 = _T_114 ? rules_57_io_n_out_12 : _GEN_1020; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1039 = _T_114 ? rules_57_io_n_out_13 : _GEN_1021; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1040 = _T_114 ? rules_57_io_n_out_14 : _GEN_1022; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1041 = _T_114 ? rules_57_io_n_out_15 : _GEN_1023; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1042 = _T_114 ? rules_57_io_n_out_16 : _GEN_1024; // @[system.scala 33:21 34:7]
  wire  _GEN_1043 = _T_114 ? rules_57_io_x_out : _GEN_1025; // @[system.scala 33:21 35:7]
  wire  _T_116 = io_en_a == 7'h3a; // @[system.scala 32:27]
  wire [1:0] _GEN_1044 = _T_116 ? rules_58_io_n_out_0 : _GEN_1026; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1045 = _T_116 ? rules_58_io_n_out_1 : _GEN_1027; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1046 = _T_116 ? rules_58_io_n_out_2 : _GEN_1028; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1047 = _T_116 ? rules_58_io_n_out_3 : _GEN_1029; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1048 = _T_116 ? rules_58_io_n_out_4 : _GEN_1030; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1049 = _T_116 ? rules_58_io_n_out_5 : _GEN_1031; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1050 = _T_116 ? rules_58_io_n_out_6 : _GEN_1032; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1051 = _T_116 ? rules_58_io_n_out_7 : _GEN_1033; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1052 = _T_116 ? rules_58_io_n_out_8 : _GEN_1034; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1053 = _T_116 ? rules_58_io_n_out_9 : _GEN_1035; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1054 = _T_116 ? rules_58_io_n_out_10 : _GEN_1036; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1055 = _T_116 ? rules_58_io_n_out_11 : _GEN_1037; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1056 = _T_116 ? rules_58_io_n_out_12 : _GEN_1038; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1057 = _T_116 ? rules_58_io_n_out_13 : _GEN_1039; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1058 = _T_116 ? rules_58_io_n_out_14 : _GEN_1040; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1059 = _T_116 ? rules_58_io_n_out_15 : _GEN_1041; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1060 = _T_116 ? rules_58_io_n_out_16 : _GEN_1042; // @[system.scala 33:21 34:7]
  wire  _GEN_1061 = _T_116 ? rules_58_io_x_out : _GEN_1043; // @[system.scala 33:21 35:7]
  wire  _T_118 = io_en_a == 7'h3b; // @[system.scala 32:27]
  wire [1:0] _GEN_1062 = _T_118 ? rules_59_io_n_out_0 : _GEN_1044; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1063 = _T_118 ? rules_59_io_n_out_1 : _GEN_1045; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1064 = _T_118 ? rules_59_io_n_out_2 : _GEN_1046; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1065 = _T_118 ? rules_59_io_n_out_3 : _GEN_1047; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1066 = _T_118 ? rules_59_io_n_out_4 : _GEN_1048; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1067 = _T_118 ? rules_59_io_n_out_5 : _GEN_1049; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1068 = _T_118 ? rules_59_io_n_out_6 : _GEN_1050; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1069 = _T_118 ? rules_59_io_n_out_7 : _GEN_1051; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1070 = _T_118 ? rules_59_io_n_out_8 : _GEN_1052; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1071 = _T_118 ? rules_59_io_n_out_9 : _GEN_1053; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1072 = _T_118 ? rules_59_io_n_out_10 : _GEN_1054; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1073 = _T_118 ? rules_59_io_n_out_11 : _GEN_1055; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1074 = _T_118 ? rules_59_io_n_out_12 : _GEN_1056; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1075 = _T_118 ? rules_59_io_n_out_13 : _GEN_1057; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1076 = _T_118 ? rules_59_io_n_out_14 : _GEN_1058; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1077 = _T_118 ? rules_59_io_n_out_15 : _GEN_1059; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1078 = _T_118 ? rules_59_io_n_out_16 : _GEN_1060; // @[system.scala 33:21 34:7]
  wire  _GEN_1079 = _T_118 ? rules_59_io_x_out : _GEN_1061; // @[system.scala 33:21 35:7]
  wire  _T_120 = io_en_a == 7'h3c; // @[system.scala 32:27]
  wire [1:0] _GEN_1080 = _T_120 ? rules_60_io_n_out_0 : _GEN_1062; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1081 = _T_120 ? rules_60_io_n_out_1 : _GEN_1063; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1082 = _T_120 ? rules_60_io_n_out_2 : _GEN_1064; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1083 = _T_120 ? rules_60_io_n_out_3 : _GEN_1065; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1084 = _T_120 ? rules_60_io_n_out_4 : _GEN_1066; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1085 = _T_120 ? rules_60_io_n_out_5 : _GEN_1067; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1086 = _T_120 ? rules_60_io_n_out_6 : _GEN_1068; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1087 = _T_120 ? rules_60_io_n_out_7 : _GEN_1069; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1088 = _T_120 ? rules_60_io_n_out_8 : _GEN_1070; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1089 = _T_120 ? rules_60_io_n_out_9 : _GEN_1071; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1090 = _T_120 ? rules_60_io_n_out_10 : _GEN_1072; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1091 = _T_120 ? rules_60_io_n_out_11 : _GEN_1073; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1092 = _T_120 ? rules_60_io_n_out_12 : _GEN_1074; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1093 = _T_120 ? rules_60_io_n_out_13 : _GEN_1075; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1094 = _T_120 ? rules_60_io_n_out_14 : _GEN_1076; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1095 = _T_120 ? rules_60_io_n_out_15 : _GEN_1077; // @[system.scala 33:21 34:7]
  wire [1:0] _GEN_1096 = _T_120 ? rules_60_io_n_out_16 : _GEN_1078; // @[system.scala 33:21 34:7]
  wire  _GEN_1097 = _T_120 ? rules_60_io_x_out : _GEN_1079; // @[system.scala 33:21 35:7]
  wire  _T_122 = io_en_a == 7'h3d; // @[system.scala 32:27]
  wire  _T_124 = io_en_a == 7'h3e; // @[system.scala 32:27]
  wire  _T_126 = io_en_a == 7'h3f; // @[system.scala 32:27]
  wire  _T_128 = io_en_a == 7'h40; // @[system.scala 32:27]
  Init rules_0 ( // @[system.scala 16:16]
    .io_en_r(rules_0_io_en_r),
    .io_n_in_0(rules_0_io_n_in_0),
    .io_n_in_1(rules_0_io_n_in_1),
    .io_n_in_2(rules_0_io_n_in_2),
    .io_n_in_3(rules_0_io_n_in_3),
    .io_n_in_4(rules_0_io_n_in_4),
    .io_n_in_5(rules_0_io_n_in_5),
    .io_n_in_6(rules_0_io_n_in_6),
    .io_n_in_7(rules_0_io_n_in_7),
    .io_n_in_8(rules_0_io_n_in_8),
    .io_n_in_9(rules_0_io_n_in_9),
    .io_n_in_10(rules_0_io_n_in_10),
    .io_n_in_11(rules_0_io_n_in_11),
    .io_n_in_12(rules_0_io_n_in_12),
    .io_n_in_13(rules_0_io_n_in_13),
    .io_n_in_14(rules_0_io_n_in_14),
    .io_n_in_15(rules_0_io_n_in_15),
    .io_n_in_16(rules_0_io_n_in_16),
    .io_n_out_0(rules_0_io_n_out_0),
    .io_n_out_1(rules_0_io_n_out_1),
    .io_n_out_2(rules_0_io_n_out_2),
    .io_n_out_3(rules_0_io_n_out_3),
    .io_n_out_4(rules_0_io_n_out_4),
    .io_n_out_5(rules_0_io_n_out_5),
    .io_n_out_6(rules_0_io_n_out_6),
    .io_n_out_7(rules_0_io_n_out_7),
    .io_n_out_8(rules_0_io_n_out_8),
    .io_n_out_9(rules_0_io_n_out_9),
    .io_n_out_10(rules_0_io_n_out_10),
    .io_n_out_11(rules_0_io_n_out_11),
    .io_n_out_12(rules_0_io_n_out_12),
    .io_n_out_13(rules_0_io_n_out_13),
    .io_n_out_14(rules_0_io_n_out_14),
    .io_n_out_15(rules_0_io_n_out_15),
    .io_n_out_16(rules_0_io_n_out_16),
    .io_x_in(rules_0_io_x_in),
    .io_x_out(rules_0_io_x_out)
  );
  Try rules_1 ( // @[system.scala 18:16]
    .io_en_r(rules_1_io_en_r),
    .io_n_in_0(rules_1_io_n_in_0),
    .io_n_in_1(rules_1_io_n_in_1),
    .io_n_in_2(rules_1_io_n_in_2),
    .io_n_in_3(rules_1_io_n_in_3),
    .io_n_in_4(rules_1_io_n_in_4),
    .io_n_in_5(rules_1_io_n_in_5),
    .io_n_in_6(rules_1_io_n_in_6),
    .io_n_in_7(rules_1_io_n_in_7),
    .io_n_in_8(rules_1_io_n_in_8),
    .io_n_in_9(rules_1_io_n_in_9),
    .io_n_in_10(rules_1_io_n_in_10),
    .io_n_in_11(rules_1_io_n_in_11),
    .io_n_in_12(rules_1_io_n_in_12),
    .io_n_in_13(rules_1_io_n_in_13),
    .io_n_in_14(rules_1_io_n_in_14),
    .io_n_in_15(rules_1_io_n_in_15),
    .io_n_in_16(rules_1_io_n_in_16),
    .io_n_out_0(rules_1_io_n_out_0),
    .io_n_out_1(rules_1_io_n_out_1),
    .io_n_out_2(rules_1_io_n_out_2),
    .io_n_out_3(rules_1_io_n_out_3),
    .io_n_out_4(rules_1_io_n_out_4),
    .io_n_out_5(rules_1_io_n_out_5),
    .io_n_out_6(rules_1_io_n_out_6),
    .io_n_out_7(rules_1_io_n_out_7),
    .io_n_out_8(rules_1_io_n_out_8),
    .io_n_out_9(rules_1_io_n_out_9),
    .io_n_out_10(rules_1_io_n_out_10),
    .io_n_out_11(rules_1_io_n_out_11),
    .io_n_out_12(rules_1_io_n_out_12),
    .io_n_out_13(rules_1_io_n_out_13),
    .io_n_out_14(rules_1_io_n_out_14),
    .io_n_out_15(rules_1_io_n_out_15),
    .io_n_out_16(rules_1_io_n_out_16),
    .io_x_in(rules_1_io_x_in),
    .io_x_out(rules_1_io_x_out)
  );
  Try_1 rules_2 ( // @[system.scala 18:16]
    .io_en_r(rules_2_io_en_r),
    .io_n_in_0(rules_2_io_n_in_0),
    .io_n_in_1(rules_2_io_n_in_1),
    .io_n_in_2(rules_2_io_n_in_2),
    .io_n_in_3(rules_2_io_n_in_3),
    .io_n_in_4(rules_2_io_n_in_4),
    .io_n_in_5(rules_2_io_n_in_5),
    .io_n_in_6(rules_2_io_n_in_6),
    .io_n_in_7(rules_2_io_n_in_7),
    .io_n_in_8(rules_2_io_n_in_8),
    .io_n_in_9(rules_2_io_n_in_9),
    .io_n_in_10(rules_2_io_n_in_10),
    .io_n_in_11(rules_2_io_n_in_11),
    .io_n_in_12(rules_2_io_n_in_12),
    .io_n_in_13(rules_2_io_n_in_13),
    .io_n_in_14(rules_2_io_n_in_14),
    .io_n_in_15(rules_2_io_n_in_15),
    .io_n_in_16(rules_2_io_n_in_16),
    .io_n_out_0(rules_2_io_n_out_0),
    .io_n_out_1(rules_2_io_n_out_1),
    .io_n_out_2(rules_2_io_n_out_2),
    .io_n_out_3(rules_2_io_n_out_3),
    .io_n_out_4(rules_2_io_n_out_4),
    .io_n_out_5(rules_2_io_n_out_5),
    .io_n_out_6(rules_2_io_n_out_6),
    .io_n_out_7(rules_2_io_n_out_7),
    .io_n_out_8(rules_2_io_n_out_8),
    .io_n_out_9(rules_2_io_n_out_9),
    .io_n_out_10(rules_2_io_n_out_10),
    .io_n_out_11(rules_2_io_n_out_11),
    .io_n_out_12(rules_2_io_n_out_12),
    .io_n_out_13(rules_2_io_n_out_13),
    .io_n_out_14(rules_2_io_n_out_14),
    .io_n_out_15(rules_2_io_n_out_15),
    .io_n_out_16(rules_2_io_n_out_16),
    .io_x_in(rules_2_io_x_in),
    .io_x_out(rules_2_io_x_out)
  );
  Try_2 rules_3 ( // @[system.scala 18:16]
    .io_en_r(rules_3_io_en_r),
    .io_n_in_0(rules_3_io_n_in_0),
    .io_n_in_1(rules_3_io_n_in_1),
    .io_n_in_2(rules_3_io_n_in_2),
    .io_n_in_3(rules_3_io_n_in_3),
    .io_n_in_4(rules_3_io_n_in_4),
    .io_n_in_5(rules_3_io_n_in_5),
    .io_n_in_6(rules_3_io_n_in_6),
    .io_n_in_7(rules_3_io_n_in_7),
    .io_n_in_8(rules_3_io_n_in_8),
    .io_n_in_9(rules_3_io_n_in_9),
    .io_n_in_10(rules_3_io_n_in_10),
    .io_n_in_11(rules_3_io_n_in_11),
    .io_n_in_12(rules_3_io_n_in_12),
    .io_n_in_13(rules_3_io_n_in_13),
    .io_n_in_14(rules_3_io_n_in_14),
    .io_n_in_15(rules_3_io_n_in_15),
    .io_n_in_16(rules_3_io_n_in_16),
    .io_n_out_0(rules_3_io_n_out_0),
    .io_n_out_1(rules_3_io_n_out_1),
    .io_n_out_2(rules_3_io_n_out_2),
    .io_n_out_3(rules_3_io_n_out_3),
    .io_n_out_4(rules_3_io_n_out_4),
    .io_n_out_5(rules_3_io_n_out_5),
    .io_n_out_6(rules_3_io_n_out_6),
    .io_n_out_7(rules_3_io_n_out_7),
    .io_n_out_8(rules_3_io_n_out_8),
    .io_n_out_9(rules_3_io_n_out_9),
    .io_n_out_10(rules_3_io_n_out_10),
    .io_n_out_11(rules_3_io_n_out_11),
    .io_n_out_12(rules_3_io_n_out_12),
    .io_n_out_13(rules_3_io_n_out_13),
    .io_n_out_14(rules_3_io_n_out_14),
    .io_n_out_15(rules_3_io_n_out_15),
    .io_n_out_16(rules_3_io_n_out_16),
    .io_x_in(rules_3_io_x_in),
    .io_x_out(rules_3_io_x_out)
  );
  Try_3 rules_4 ( // @[system.scala 18:16]
    .io_en_r(rules_4_io_en_r),
    .io_n_in_0(rules_4_io_n_in_0),
    .io_n_in_1(rules_4_io_n_in_1),
    .io_n_in_2(rules_4_io_n_in_2),
    .io_n_in_3(rules_4_io_n_in_3),
    .io_n_in_4(rules_4_io_n_in_4),
    .io_n_in_5(rules_4_io_n_in_5),
    .io_n_in_6(rules_4_io_n_in_6),
    .io_n_in_7(rules_4_io_n_in_7),
    .io_n_in_8(rules_4_io_n_in_8),
    .io_n_in_9(rules_4_io_n_in_9),
    .io_n_in_10(rules_4_io_n_in_10),
    .io_n_in_11(rules_4_io_n_in_11),
    .io_n_in_12(rules_4_io_n_in_12),
    .io_n_in_13(rules_4_io_n_in_13),
    .io_n_in_14(rules_4_io_n_in_14),
    .io_n_in_15(rules_4_io_n_in_15),
    .io_n_in_16(rules_4_io_n_in_16),
    .io_n_out_0(rules_4_io_n_out_0),
    .io_n_out_1(rules_4_io_n_out_1),
    .io_n_out_2(rules_4_io_n_out_2),
    .io_n_out_3(rules_4_io_n_out_3),
    .io_n_out_4(rules_4_io_n_out_4),
    .io_n_out_5(rules_4_io_n_out_5),
    .io_n_out_6(rules_4_io_n_out_6),
    .io_n_out_7(rules_4_io_n_out_7),
    .io_n_out_8(rules_4_io_n_out_8),
    .io_n_out_9(rules_4_io_n_out_9),
    .io_n_out_10(rules_4_io_n_out_10),
    .io_n_out_11(rules_4_io_n_out_11),
    .io_n_out_12(rules_4_io_n_out_12),
    .io_n_out_13(rules_4_io_n_out_13),
    .io_n_out_14(rules_4_io_n_out_14),
    .io_n_out_15(rules_4_io_n_out_15),
    .io_n_out_16(rules_4_io_n_out_16),
    .io_x_in(rules_4_io_x_in),
    .io_x_out(rules_4_io_x_out)
  );
  Try_4 rules_5 ( // @[system.scala 18:16]
    .io_en_r(rules_5_io_en_r),
    .io_n_in_0(rules_5_io_n_in_0),
    .io_n_in_1(rules_5_io_n_in_1),
    .io_n_in_2(rules_5_io_n_in_2),
    .io_n_in_3(rules_5_io_n_in_3),
    .io_n_in_4(rules_5_io_n_in_4),
    .io_n_in_5(rules_5_io_n_in_5),
    .io_n_in_6(rules_5_io_n_in_6),
    .io_n_in_7(rules_5_io_n_in_7),
    .io_n_in_8(rules_5_io_n_in_8),
    .io_n_in_9(rules_5_io_n_in_9),
    .io_n_in_10(rules_5_io_n_in_10),
    .io_n_in_11(rules_5_io_n_in_11),
    .io_n_in_12(rules_5_io_n_in_12),
    .io_n_in_13(rules_5_io_n_in_13),
    .io_n_in_14(rules_5_io_n_in_14),
    .io_n_in_15(rules_5_io_n_in_15),
    .io_n_in_16(rules_5_io_n_in_16),
    .io_n_out_0(rules_5_io_n_out_0),
    .io_n_out_1(rules_5_io_n_out_1),
    .io_n_out_2(rules_5_io_n_out_2),
    .io_n_out_3(rules_5_io_n_out_3),
    .io_n_out_4(rules_5_io_n_out_4),
    .io_n_out_5(rules_5_io_n_out_5),
    .io_n_out_6(rules_5_io_n_out_6),
    .io_n_out_7(rules_5_io_n_out_7),
    .io_n_out_8(rules_5_io_n_out_8),
    .io_n_out_9(rules_5_io_n_out_9),
    .io_n_out_10(rules_5_io_n_out_10),
    .io_n_out_11(rules_5_io_n_out_11),
    .io_n_out_12(rules_5_io_n_out_12),
    .io_n_out_13(rules_5_io_n_out_13),
    .io_n_out_14(rules_5_io_n_out_14),
    .io_n_out_15(rules_5_io_n_out_15),
    .io_n_out_16(rules_5_io_n_out_16),
    .io_x_in(rules_5_io_x_in),
    .io_x_out(rules_5_io_x_out)
  );
  Try_5 rules_6 ( // @[system.scala 18:16]
    .io_en_r(rules_6_io_en_r),
    .io_n_in_0(rules_6_io_n_in_0),
    .io_n_in_1(rules_6_io_n_in_1),
    .io_n_in_2(rules_6_io_n_in_2),
    .io_n_in_3(rules_6_io_n_in_3),
    .io_n_in_4(rules_6_io_n_in_4),
    .io_n_in_5(rules_6_io_n_in_5),
    .io_n_in_6(rules_6_io_n_in_6),
    .io_n_in_7(rules_6_io_n_in_7),
    .io_n_in_8(rules_6_io_n_in_8),
    .io_n_in_9(rules_6_io_n_in_9),
    .io_n_in_10(rules_6_io_n_in_10),
    .io_n_in_11(rules_6_io_n_in_11),
    .io_n_in_12(rules_6_io_n_in_12),
    .io_n_in_13(rules_6_io_n_in_13),
    .io_n_in_14(rules_6_io_n_in_14),
    .io_n_in_15(rules_6_io_n_in_15),
    .io_n_in_16(rules_6_io_n_in_16),
    .io_n_out_0(rules_6_io_n_out_0),
    .io_n_out_1(rules_6_io_n_out_1),
    .io_n_out_2(rules_6_io_n_out_2),
    .io_n_out_3(rules_6_io_n_out_3),
    .io_n_out_4(rules_6_io_n_out_4),
    .io_n_out_5(rules_6_io_n_out_5),
    .io_n_out_6(rules_6_io_n_out_6),
    .io_n_out_7(rules_6_io_n_out_7),
    .io_n_out_8(rules_6_io_n_out_8),
    .io_n_out_9(rules_6_io_n_out_9),
    .io_n_out_10(rules_6_io_n_out_10),
    .io_n_out_11(rules_6_io_n_out_11),
    .io_n_out_12(rules_6_io_n_out_12),
    .io_n_out_13(rules_6_io_n_out_13),
    .io_n_out_14(rules_6_io_n_out_14),
    .io_n_out_15(rules_6_io_n_out_15),
    .io_n_out_16(rules_6_io_n_out_16),
    .io_x_in(rules_6_io_x_in),
    .io_x_out(rules_6_io_x_out)
  );
  Try_6 rules_7 ( // @[system.scala 18:16]
    .io_en_r(rules_7_io_en_r),
    .io_n_in_0(rules_7_io_n_in_0),
    .io_n_in_1(rules_7_io_n_in_1),
    .io_n_in_2(rules_7_io_n_in_2),
    .io_n_in_3(rules_7_io_n_in_3),
    .io_n_in_4(rules_7_io_n_in_4),
    .io_n_in_5(rules_7_io_n_in_5),
    .io_n_in_6(rules_7_io_n_in_6),
    .io_n_in_7(rules_7_io_n_in_7),
    .io_n_in_8(rules_7_io_n_in_8),
    .io_n_in_9(rules_7_io_n_in_9),
    .io_n_in_10(rules_7_io_n_in_10),
    .io_n_in_11(rules_7_io_n_in_11),
    .io_n_in_12(rules_7_io_n_in_12),
    .io_n_in_13(rules_7_io_n_in_13),
    .io_n_in_14(rules_7_io_n_in_14),
    .io_n_in_15(rules_7_io_n_in_15),
    .io_n_in_16(rules_7_io_n_in_16),
    .io_n_out_0(rules_7_io_n_out_0),
    .io_n_out_1(rules_7_io_n_out_1),
    .io_n_out_2(rules_7_io_n_out_2),
    .io_n_out_3(rules_7_io_n_out_3),
    .io_n_out_4(rules_7_io_n_out_4),
    .io_n_out_5(rules_7_io_n_out_5),
    .io_n_out_6(rules_7_io_n_out_6),
    .io_n_out_7(rules_7_io_n_out_7),
    .io_n_out_8(rules_7_io_n_out_8),
    .io_n_out_9(rules_7_io_n_out_9),
    .io_n_out_10(rules_7_io_n_out_10),
    .io_n_out_11(rules_7_io_n_out_11),
    .io_n_out_12(rules_7_io_n_out_12),
    .io_n_out_13(rules_7_io_n_out_13),
    .io_n_out_14(rules_7_io_n_out_14),
    .io_n_out_15(rules_7_io_n_out_15),
    .io_n_out_16(rules_7_io_n_out_16),
    .io_x_in(rules_7_io_x_in),
    .io_x_out(rules_7_io_x_out)
  );
  Try_7 rules_8 ( // @[system.scala 18:16]
    .io_en_r(rules_8_io_en_r),
    .io_n_in_0(rules_8_io_n_in_0),
    .io_n_in_1(rules_8_io_n_in_1),
    .io_n_in_2(rules_8_io_n_in_2),
    .io_n_in_3(rules_8_io_n_in_3),
    .io_n_in_4(rules_8_io_n_in_4),
    .io_n_in_5(rules_8_io_n_in_5),
    .io_n_in_6(rules_8_io_n_in_6),
    .io_n_in_7(rules_8_io_n_in_7),
    .io_n_in_8(rules_8_io_n_in_8),
    .io_n_in_9(rules_8_io_n_in_9),
    .io_n_in_10(rules_8_io_n_in_10),
    .io_n_in_11(rules_8_io_n_in_11),
    .io_n_in_12(rules_8_io_n_in_12),
    .io_n_in_13(rules_8_io_n_in_13),
    .io_n_in_14(rules_8_io_n_in_14),
    .io_n_in_15(rules_8_io_n_in_15),
    .io_n_in_16(rules_8_io_n_in_16),
    .io_n_out_0(rules_8_io_n_out_0),
    .io_n_out_1(rules_8_io_n_out_1),
    .io_n_out_2(rules_8_io_n_out_2),
    .io_n_out_3(rules_8_io_n_out_3),
    .io_n_out_4(rules_8_io_n_out_4),
    .io_n_out_5(rules_8_io_n_out_5),
    .io_n_out_6(rules_8_io_n_out_6),
    .io_n_out_7(rules_8_io_n_out_7),
    .io_n_out_8(rules_8_io_n_out_8),
    .io_n_out_9(rules_8_io_n_out_9),
    .io_n_out_10(rules_8_io_n_out_10),
    .io_n_out_11(rules_8_io_n_out_11),
    .io_n_out_12(rules_8_io_n_out_12),
    .io_n_out_13(rules_8_io_n_out_13),
    .io_n_out_14(rules_8_io_n_out_14),
    .io_n_out_15(rules_8_io_n_out_15),
    .io_n_out_16(rules_8_io_n_out_16),
    .io_x_in(rules_8_io_x_in),
    .io_x_out(rules_8_io_x_out)
  );
  Try_8 rules_9 ( // @[system.scala 18:16]
    .io_en_r(rules_9_io_en_r),
    .io_n_in_0(rules_9_io_n_in_0),
    .io_n_in_1(rules_9_io_n_in_1),
    .io_n_in_2(rules_9_io_n_in_2),
    .io_n_in_3(rules_9_io_n_in_3),
    .io_n_in_4(rules_9_io_n_in_4),
    .io_n_in_5(rules_9_io_n_in_5),
    .io_n_in_6(rules_9_io_n_in_6),
    .io_n_in_7(rules_9_io_n_in_7),
    .io_n_in_8(rules_9_io_n_in_8),
    .io_n_in_9(rules_9_io_n_in_9),
    .io_n_in_10(rules_9_io_n_in_10),
    .io_n_in_11(rules_9_io_n_in_11),
    .io_n_in_12(rules_9_io_n_in_12),
    .io_n_in_13(rules_9_io_n_in_13),
    .io_n_in_14(rules_9_io_n_in_14),
    .io_n_in_15(rules_9_io_n_in_15),
    .io_n_in_16(rules_9_io_n_in_16),
    .io_n_out_0(rules_9_io_n_out_0),
    .io_n_out_1(rules_9_io_n_out_1),
    .io_n_out_2(rules_9_io_n_out_2),
    .io_n_out_3(rules_9_io_n_out_3),
    .io_n_out_4(rules_9_io_n_out_4),
    .io_n_out_5(rules_9_io_n_out_5),
    .io_n_out_6(rules_9_io_n_out_6),
    .io_n_out_7(rules_9_io_n_out_7),
    .io_n_out_8(rules_9_io_n_out_8),
    .io_n_out_9(rules_9_io_n_out_9),
    .io_n_out_10(rules_9_io_n_out_10),
    .io_n_out_11(rules_9_io_n_out_11),
    .io_n_out_12(rules_9_io_n_out_12),
    .io_n_out_13(rules_9_io_n_out_13),
    .io_n_out_14(rules_9_io_n_out_14),
    .io_n_out_15(rules_9_io_n_out_15),
    .io_n_out_16(rules_9_io_n_out_16),
    .io_x_in(rules_9_io_x_in),
    .io_x_out(rules_9_io_x_out)
  );
  Try_9 rules_10 ( // @[system.scala 18:16]
    .io_en_r(rules_10_io_en_r),
    .io_n_in_0(rules_10_io_n_in_0),
    .io_n_in_1(rules_10_io_n_in_1),
    .io_n_in_2(rules_10_io_n_in_2),
    .io_n_in_3(rules_10_io_n_in_3),
    .io_n_in_4(rules_10_io_n_in_4),
    .io_n_in_5(rules_10_io_n_in_5),
    .io_n_in_6(rules_10_io_n_in_6),
    .io_n_in_7(rules_10_io_n_in_7),
    .io_n_in_8(rules_10_io_n_in_8),
    .io_n_in_9(rules_10_io_n_in_9),
    .io_n_in_10(rules_10_io_n_in_10),
    .io_n_in_11(rules_10_io_n_in_11),
    .io_n_in_12(rules_10_io_n_in_12),
    .io_n_in_13(rules_10_io_n_in_13),
    .io_n_in_14(rules_10_io_n_in_14),
    .io_n_in_15(rules_10_io_n_in_15),
    .io_n_in_16(rules_10_io_n_in_16),
    .io_n_out_0(rules_10_io_n_out_0),
    .io_n_out_1(rules_10_io_n_out_1),
    .io_n_out_2(rules_10_io_n_out_2),
    .io_n_out_3(rules_10_io_n_out_3),
    .io_n_out_4(rules_10_io_n_out_4),
    .io_n_out_5(rules_10_io_n_out_5),
    .io_n_out_6(rules_10_io_n_out_6),
    .io_n_out_7(rules_10_io_n_out_7),
    .io_n_out_8(rules_10_io_n_out_8),
    .io_n_out_9(rules_10_io_n_out_9),
    .io_n_out_10(rules_10_io_n_out_10),
    .io_n_out_11(rules_10_io_n_out_11),
    .io_n_out_12(rules_10_io_n_out_12),
    .io_n_out_13(rules_10_io_n_out_13),
    .io_n_out_14(rules_10_io_n_out_14),
    .io_n_out_15(rules_10_io_n_out_15),
    .io_n_out_16(rules_10_io_n_out_16),
    .io_x_in(rules_10_io_x_in),
    .io_x_out(rules_10_io_x_out)
  );
  Try_10 rules_11 ( // @[system.scala 18:16]
    .io_en_r(rules_11_io_en_r),
    .io_n_in_0(rules_11_io_n_in_0),
    .io_n_in_1(rules_11_io_n_in_1),
    .io_n_in_2(rules_11_io_n_in_2),
    .io_n_in_3(rules_11_io_n_in_3),
    .io_n_in_4(rules_11_io_n_in_4),
    .io_n_in_5(rules_11_io_n_in_5),
    .io_n_in_6(rules_11_io_n_in_6),
    .io_n_in_7(rules_11_io_n_in_7),
    .io_n_in_8(rules_11_io_n_in_8),
    .io_n_in_9(rules_11_io_n_in_9),
    .io_n_in_10(rules_11_io_n_in_10),
    .io_n_in_11(rules_11_io_n_in_11),
    .io_n_in_12(rules_11_io_n_in_12),
    .io_n_in_13(rules_11_io_n_in_13),
    .io_n_in_14(rules_11_io_n_in_14),
    .io_n_in_15(rules_11_io_n_in_15),
    .io_n_in_16(rules_11_io_n_in_16),
    .io_n_out_0(rules_11_io_n_out_0),
    .io_n_out_1(rules_11_io_n_out_1),
    .io_n_out_2(rules_11_io_n_out_2),
    .io_n_out_3(rules_11_io_n_out_3),
    .io_n_out_4(rules_11_io_n_out_4),
    .io_n_out_5(rules_11_io_n_out_5),
    .io_n_out_6(rules_11_io_n_out_6),
    .io_n_out_7(rules_11_io_n_out_7),
    .io_n_out_8(rules_11_io_n_out_8),
    .io_n_out_9(rules_11_io_n_out_9),
    .io_n_out_10(rules_11_io_n_out_10),
    .io_n_out_11(rules_11_io_n_out_11),
    .io_n_out_12(rules_11_io_n_out_12),
    .io_n_out_13(rules_11_io_n_out_13),
    .io_n_out_14(rules_11_io_n_out_14),
    .io_n_out_15(rules_11_io_n_out_15),
    .io_n_out_16(rules_11_io_n_out_16),
    .io_x_in(rules_11_io_x_in),
    .io_x_out(rules_11_io_x_out)
  );
  Try_11 rules_12 ( // @[system.scala 18:16]
    .io_en_r(rules_12_io_en_r),
    .io_n_in_0(rules_12_io_n_in_0),
    .io_n_in_1(rules_12_io_n_in_1),
    .io_n_in_2(rules_12_io_n_in_2),
    .io_n_in_3(rules_12_io_n_in_3),
    .io_n_in_4(rules_12_io_n_in_4),
    .io_n_in_5(rules_12_io_n_in_5),
    .io_n_in_6(rules_12_io_n_in_6),
    .io_n_in_7(rules_12_io_n_in_7),
    .io_n_in_8(rules_12_io_n_in_8),
    .io_n_in_9(rules_12_io_n_in_9),
    .io_n_in_10(rules_12_io_n_in_10),
    .io_n_in_11(rules_12_io_n_in_11),
    .io_n_in_12(rules_12_io_n_in_12),
    .io_n_in_13(rules_12_io_n_in_13),
    .io_n_in_14(rules_12_io_n_in_14),
    .io_n_in_15(rules_12_io_n_in_15),
    .io_n_in_16(rules_12_io_n_in_16),
    .io_n_out_0(rules_12_io_n_out_0),
    .io_n_out_1(rules_12_io_n_out_1),
    .io_n_out_2(rules_12_io_n_out_2),
    .io_n_out_3(rules_12_io_n_out_3),
    .io_n_out_4(rules_12_io_n_out_4),
    .io_n_out_5(rules_12_io_n_out_5),
    .io_n_out_6(rules_12_io_n_out_6),
    .io_n_out_7(rules_12_io_n_out_7),
    .io_n_out_8(rules_12_io_n_out_8),
    .io_n_out_9(rules_12_io_n_out_9),
    .io_n_out_10(rules_12_io_n_out_10),
    .io_n_out_11(rules_12_io_n_out_11),
    .io_n_out_12(rules_12_io_n_out_12),
    .io_n_out_13(rules_12_io_n_out_13),
    .io_n_out_14(rules_12_io_n_out_14),
    .io_n_out_15(rules_12_io_n_out_15),
    .io_n_out_16(rules_12_io_n_out_16),
    .io_x_in(rules_12_io_x_in),
    .io_x_out(rules_12_io_x_out)
  );
  Try_12 rules_13 ( // @[system.scala 18:16]
    .io_en_r(rules_13_io_en_r),
    .io_n_in_0(rules_13_io_n_in_0),
    .io_n_in_1(rules_13_io_n_in_1),
    .io_n_in_2(rules_13_io_n_in_2),
    .io_n_in_3(rules_13_io_n_in_3),
    .io_n_in_4(rules_13_io_n_in_4),
    .io_n_in_5(rules_13_io_n_in_5),
    .io_n_in_6(rules_13_io_n_in_6),
    .io_n_in_7(rules_13_io_n_in_7),
    .io_n_in_8(rules_13_io_n_in_8),
    .io_n_in_9(rules_13_io_n_in_9),
    .io_n_in_10(rules_13_io_n_in_10),
    .io_n_in_11(rules_13_io_n_in_11),
    .io_n_in_12(rules_13_io_n_in_12),
    .io_n_in_13(rules_13_io_n_in_13),
    .io_n_in_14(rules_13_io_n_in_14),
    .io_n_in_15(rules_13_io_n_in_15),
    .io_n_in_16(rules_13_io_n_in_16),
    .io_n_out_0(rules_13_io_n_out_0),
    .io_n_out_1(rules_13_io_n_out_1),
    .io_n_out_2(rules_13_io_n_out_2),
    .io_n_out_3(rules_13_io_n_out_3),
    .io_n_out_4(rules_13_io_n_out_4),
    .io_n_out_5(rules_13_io_n_out_5),
    .io_n_out_6(rules_13_io_n_out_6),
    .io_n_out_7(rules_13_io_n_out_7),
    .io_n_out_8(rules_13_io_n_out_8),
    .io_n_out_9(rules_13_io_n_out_9),
    .io_n_out_10(rules_13_io_n_out_10),
    .io_n_out_11(rules_13_io_n_out_11),
    .io_n_out_12(rules_13_io_n_out_12),
    .io_n_out_13(rules_13_io_n_out_13),
    .io_n_out_14(rules_13_io_n_out_14),
    .io_n_out_15(rules_13_io_n_out_15),
    .io_n_out_16(rules_13_io_n_out_16),
    .io_x_in(rules_13_io_x_in),
    .io_x_out(rules_13_io_x_out)
  );
  Try_13 rules_14 ( // @[system.scala 18:16]
    .io_en_r(rules_14_io_en_r),
    .io_n_in_0(rules_14_io_n_in_0),
    .io_n_in_1(rules_14_io_n_in_1),
    .io_n_in_2(rules_14_io_n_in_2),
    .io_n_in_3(rules_14_io_n_in_3),
    .io_n_in_4(rules_14_io_n_in_4),
    .io_n_in_5(rules_14_io_n_in_5),
    .io_n_in_6(rules_14_io_n_in_6),
    .io_n_in_7(rules_14_io_n_in_7),
    .io_n_in_8(rules_14_io_n_in_8),
    .io_n_in_9(rules_14_io_n_in_9),
    .io_n_in_10(rules_14_io_n_in_10),
    .io_n_in_11(rules_14_io_n_in_11),
    .io_n_in_12(rules_14_io_n_in_12),
    .io_n_in_13(rules_14_io_n_in_13),
    .io_n_in_14(rules_14_io_n_in_14),
    .io_n_in_15(rules_14_io_n_in_15),
    .io_n_in_16(rules_14_io_n_in_16),
    .io_n_out_0(rules_14_io_n_out_0),
    .io_n_out_1(rules_14_io_n_out_1),
    .io_n_out_2(rules_14_io_n_out_2),
    .io_n_out_3(rules_14_io_n_out_3),
    .io_n_out_4(rules_14_io_n_out_4),
    .io_n_out_5(rules_14_io_n_out_5),
    .io_n_out_6(rules_14_io_n_out_6),
    .io_n_out_7(rules_14_io_n_out_7),
    .io_n_out_8(rules_14_io_n_out_8),
    .io_n_out_9(rules_14_io_n_out_9),
    .io_n_out_10(rules_14_io_n_out_10),
    .io_n_out_11(rules_14_io_n_out_11),
    .io_n_out_12(rules_14_io_n_out_12),
    .io_n_out_13(rules_14_io_n_out_13),
    .io_n_out_14(rules_14_io_n_out_14),
    .io_n_out_15(rules_14_io_n_out_15),
    .io_n_out_16(rules_14_io_n_out_16),
    .io_x_in(rules_14_io_x_in),
    .io_x_out(rules_14_io_x_out)
  );
  Try_14 rules_15 ( // @[system.scala 18:16]
    .io_en_r(rules_15_io_en_r),
    .io_n_in_0(rules_15_io_n_in_0),
    .io_n_in_1(rules_15_io_n_in_1),
    .io_n_in_2(rules_15_io_n_in_2),
    .io_n_in_3(rules_15_io_n_in_3),
    .io_n_in_4(rules_15_io_n_in_4),
    .io_n_in_5(rules_15_io_n_in_5),
    .io_n_in_6(rules_15_io_n_in_6),
    .io_n_in_7(rules_15_io_n_in_7),
    .io_n_in_8(rules_15_io_n_in_8),
    .io_n_in_9(rules_15_io_n_in_9),
    .io_n_in_10(rules_15_io_n_in_10),
    .io_n_in_11(rules_15_io_n_in_11),
    .io_n_in_12(rules_15_io_n_in_12),
    .io_n_in_13(rules_15_io_n_in_13),
    .io_n_in_14(rules_15_io_n_in_14),
    .io_n_in_15(rules_15_io_n_in_15),
    .io_n_in_16(rules_15_io_n_in_16),
    .io_n_out_0(rules_15_io_n_out_0),
    .io_n_out_1(rules_15_io_n_out_1),
    .io_n_out_2(rules_15_io_n_out_2),
    .io_n_out_3(rules_15_io_n_out_3),
    .io_n_out_4(rules_15_io_n_out_4),
    .io_n_out_5(rules_15_io_n_out_5),
    .io_n_out_6(rules_15_io_n_out_6),
    .io_n_out_7(rules_15_io_n_out_7),
    .io_n_out_8(rules_15_io_n_out_8),
    .io_n_out_9(rules_15_io_n_out_9),
    .io_n_out_10(rules_15_io_n_out_10),
    .io_n_out_11(rules_15_io_n_out_11),
    .io_n_out_12(rules_15_io_n_out_12),
    .io_n_out_13(rules_15_io_n_out_13),
    .io_n_out_14(rules_15_io_n_out_14),
    .io_n_out_15(rules_15_io_n_out_15),
    .io_n_out_16(rules_15_io_n_out_16),
    .io_x_in(rules_15_io_x_in),
    .io_x_out(rules_15_io_x_out)
  );
  Try_15 rules_16 ( // @[system.scala 18:16]
    .io_en_r(rules_16_io_en_r),
    .io_n_in_0(rules_16_io_n_in_0),
    .io_n_in_1(rules_16_io_n_in_1),
    .io_n_in_2(rules_16_io_n_in_2),
    .io_n_in_3(rules_16_io_n_in_3),
    .io_n_in_4(rules_16_io_n_in_4),
    .io_n_in_5(rules_16_io_n_in_5),
    .io_n_in_6(rules_16_io_n_in_6),
    .io_n_in_7(rules_16_io_n_in_7),
    .io_n_in_8(rules_16_io_n_in_8),
    .io_n_in_9(rules_16_io_n_in_9),
    .io_n_in_10(rules_16_io_n_in_10),
    .io_n_in_11(rules_16_io_n_in_11),
    .io_n_in_12(rules_16_io_n_in_12),
    .io_n_in_13(rules_16_io_n_in_13),
    .io_n_in_14(rules_16_io_n_in_14),
    .io_n_in_15(rules_16_io_n_in_15),
    .io_n_in_16(rules_16_io_n_in_16),
    .io_n_out_0(rules_16_io_n_out_0),
    .io_n_out_1(rules_16_io_n_out_1),
    .io_n_out_2(rules_16_io_n_out_2),
    .io_n_out_3(rules_16_io_n_out_3),
    .io_n_out_4(rules_16_io_n_out_4),
    .io_n_out_5(rules_16_io_n_out_5),
    .io_n_out_6(rules_16_io_n_out_6),
    .io_n_out_7(rules_16_io_n_out_7),
    .io_n_out_8(rules_16_io_n_out_8),
    .io_n_out_9(rules_16_io_n_out_9),
    .io_n_out_10(rules_16_io_n_out_10),
    .io_n_out_11(rules_16_io_n_out_11),
    .io_n_out_12(rules_16_io_n_out_12),
    .io_n_out_13(rules_16_io_n_out_13),
    .io_n_out_14(rules_16_io_n_out_14),
    .io_n_out_15(rules_16_io_n_out_15),
    .io_n_out_16(rules_16_io_n_out_16),
    .io_x_in(rules_16_io_x_in),
    .io_x_out(rules_16_io_x_out)
  );
  Crit rules_17 ( // @[system.scala 21:16]
    .io_en_r(rules_17_io_en_r),
    .io_n_in_0(rules_17_io_n_in_0),
    .io_n_in_1(rules_17_io_n_in_1),
    .io_n_in_2(rules_17_io_n_in_2),
    .io_n_in_3(rules_17_io_n_in_3),
    .io_n_in_4(rules_17_io_n_in_4),
    .io_n_in_5(rules_17_io_n_in_5),
    .io_n_in_6(rules_17_io_n_in_6),
    .io_n_in_7(rules_17_io_n_in_7),
    .io_n_in_8(rules_17_io_n_in_8),
    .io_n_in_9(rules_17_io_n_in_9),
    .io_n_in_10(rules_17_io_n_in_10),
    .io_n_in_11(rules_17_io_n_in_11),
    .io_n_in_12(rules_17_io_n_in_12),
    .io_n_in_13(rules_17_io_n_in_13),
    .io_n_in_14(rules_17_io_n_in_14),
    .io_n_in_15(rules_17_io_n_in_15),
    .io_n_in_16(rules_17_io_n_in_16),
    .io_n_out_0(rules_17_io_n_out_0),
    .io_n_out_1(rules_17_io_n_out_1),
    .io_n_out_2(rules_17_io_n_out_2),
    .io_n_out_3(rules_17_io_n_out_3),
    .io_n_out_4(rules_17_io_n_out_4),
    .io_n_out_5(rules_17_io_n_out_5),
    .io_n_out_6(rules_17_io_n_out_6),
    .io_n_out_7(rules_17_io_n_out_7),
    .io_n_out_8(rules_17_io_n_out_8),
    .io_n_out_9(rules_17_io_n_out_9),
    .io_n_out_10(rules_17_io_n_out_10),
    .io_n_out_11(rules_17_io_n_out_11),
    .io_n_out_12(rules_17_io_n_out_12),
    .io_n_out_13(rules_17_io_n_out_13),
    .io_n_out_14(rules_17_io_n_out_14),
    .io_n_out_15(rules_17_io_n_out_15),
    .io_n_out_16(rules_17_io_n_out_16),
    .io_x_in(rules_17_io_x_in),
    .io_x_out(rules_17_io_x_out)
  );
  Crit_1 rules_18 ( // @[system.scala 21:16]
    .io_en_r(rules_18_io_en_r),
    .io_n_in_0(rules_18_io_n_in_0),
    .io_n_in_1(rules_18_io_n_in_1),
    .io_n_in_2(rules_18_io_n_in_2),
    .io_n_in_3(rules_18_io_n_in_3),
    .io_n_in_4(rules_18_io_n_in_4),
    .io_n_in_5(rules_18_io_n_in_5),
    .io_n_in_6(rules_18_io_n_in_6),
    .io_n_in_7(rules_18_io_n_in_7),
    .io_n_in_8(rules_18_io_n_in_8),
    .io_n_in_9(rules_18_io_n_in_9),
    .io_n_in_10(rules_18_io_n_in_10),
    .io_n_in_11(rules_18_io_n_in_11),
    .io_n_in_12(rules_18_io_n_in_12),
    .io_n_in_13(rules_18_io_n_in_13),
    .io_n_in_14(rules_18_io_n_in_14),
    .io_n_in_15(rules_18_io_n_in_15),
    .io_n_in_16(rules_18_io_n_in_16),
    .io_n_out_0(rules_18_io_n_out_0),
    .io_n_out_1(rules_18_io_n_out_1),
    .io_n_out_2(rules_18_io_n_out_2),
    .io_n_out_3(rules_18_io_n_out_3),
    .io_n_out_4(rules_18_io_n_out_4),
    .io_n_out_5(rules_18_io_n_out_5),
    .io_n_out_6(rules_18_io_n_out_6),
    .io_n_out_7(rules_18_io_n_out_7),
    .io_n_out_8(rules_18_io_n_out_8),
    .io_n_out_9(rules_18_io_n_out_9),
    .io_n_out_10(rules_18_io_n_out_10),
    .io_n_out_11(rules_18_io_n_out_11),
    .io_n_out_12(rules_18_io_n_out_12),
    .io_n_out_13(rules_18_io_n_out_13),
    .io_n_out_14(rules_18_io_n_out_14),
    .io_n_out_15(rules_18_io_n_out_15),
    .io_n_out_16(rules_18_io_n_out_16),
    .io_x_in(rules_18_io_x_in),
    .io_x_out(rules_18_io_x_out)
  );
  Crit_2 rules_19 ( // @[system.scala 21:16]
    .io_en_r(rules_19_io_en_r),
    .io_n_in_0(rules_19_io_n_in_0),
    .io_n_in_1(rules_19_io_n_in_1),
    .io_n_in_2(rules_19_io_n_in_2),
    .io_n_in_3(rules_19_io_n_in_3),
    .io_n_in_4(rules_19_io_n_in_4),
    .io_n_in_5(rules_19_io_n_in_5),
    .io_n_in_6(rules_19_io_n_in_6),
    .io_n_in_7(rules_19_io_n_in_7),
    .io_n_in_8(rules_19_io_n_in_8),
    .io_n_in_9(rules_19_io_n_in_9),
    .io_n_in_10(rules_19_io_n_in_10),
    .io_n_in_11(rules_19_io_n_in_11),
    .io_n_in_12(rules_19_io_n_in_12),
    .io_n_in_13(rules_19_io_n_in_13),
    .io_n_in_14(rules_19_io_n_in_14),
    .io_n_in_15(rules_19_io_n_in_15),
    .io_n_in_16(rules_19_io_n_in_16),
    .io_n_out_0(rules_19_io_n_out_0),
    .io_n_out_1(rules_19_io_n_out_1),
    .io_n_out_2(rules_19_io_n_out_2),
    .io_n_out_3(rules_19_io_n_out_3),
    .io_n_out_4(rules_19_io_n_out_4),
    .io_n_out_5(rules_19_io_n_out_5),
    .io_n_out_6(rules_19_io_n_out_6),
    .io_n_out_7(rules_19_io_n_out_7),
    .io_n_out_8(rules_19_io_n_out_8),
    .io_n_out_9(rules_19_io_n_out_9),
    .io_n_out_10(rules_19_io_n_out_10),
    .io_n_out_11(rules_19_io_n_out_11),
    .io_n_out_12(rules_19_io_n_out_12),
    .io_n_out_13(rules_19_io_n_out_13),
    .io_n_out_14(rules_19_io_n_out_14),
    .io_n_out_15(rules_19_io_n_out_15),
    .io_n_out_16(rules_19_io_n_out_16),
    .io_x_in(rules_19_io_x_in),
    .io_x_out(rules_19_io_x_out)
  );
  Crit_3 rules_20 ( // @[system.scala 21:16]
    .io_en_r(rules_20_io_en_r),
    .io_n_in_0(rules_20_io_n_in_0),
    .io_n_in_1(rules_20_io_n_in_1),
    .io_n_in_2(rules_20_io_n_in_2),
    .io_n_in_3(rules_20_io_n_in_3),
    .io_n_in_4(rules_20_io_n_in_4),
    .io_n_in_5(rules_20_io_n_in_5),
    .io_n_in_6(rules_20_io_n_in_6),
    .io_n_in_7(rules_20_io_n_in_7),
    .io_n_in_8(rules_20_io_n_in_8),
    .io_n_in_9(rules_20_io_n_in_9),
    .io_n_in_10(rules_20_io_n_in_10),
    .io_n_in_11(rules_20_io_n_in_11),
    .io_n_in_12(rules_20_io_n_in_12),
    .io_n_in_13(rules_20_io_n_in_13),
    .io_n_in_14(rules_20_io_n_in_14),
    .io_n_in_15(rules_20_io_n_in_15),
    .io_n_in_16(rules_20_io_n_in_16),
    .io_n_out_0(rules_20_io_n_out_0),
    .io_n_out_1(rules_20_io_n_out_1),
    .io_n_out_2(rules_20_io_n_out_2),
    .io_n_out_3(rules_20_io_n_out_3),
    .io_n_out_4(rules_20_io_n_out_4),
    .io_n_out_5(rules_20_io_n_out_5),
    .io_n_out_6(rules_20_io_n_out_6),
    .io_n_out_7(rules_20_io_n_out_7),
    .io_n_out_8(rules_20_io_n_out_8),
    .io_n_out_9(rules_20_io_n_out_9),
    .io_n_out_10(rules_20_io_n_out_10),
    .io_n_out_11(rules_20_io_n_out_11),
    .io_n_out_12(rules_20_io_n_out_12),
    .io_n_out_13(rules_20_io_n_out_13),
    .io_n_out_14(rules_20_io_n_out_14),
    .io_n_out_15(rules_20_io_n_out_15),
    .io_n_out_16(rules_20_io_n_out_16),
    .io_x_in(rules_20_io_x_in),
    .io_x_out(rules_20_io_x_out)
  );
  Crit_4 rules_21 ( // @[system.scala 21:16]
    .io_en_r(rules_21_io_en_r),
    .io_n_in_0(rules_21_io_n_in_0),
    .io_n_in_1(rules_21_io_n_in_1),
    .io_n_in_2(rules_21_io_n_in_2),
    .io_n_in_3(rules_21_io_n_in_3),
    .io_n_in_4(rules_21_io_n_in_4),
    .io_n_in_5(rules_21_io_n_in_5),
    .io_n_in_6(rules_21_io_n_in_6),
    .io_n_in_7(rules_21_io_n_in_7),
    .io_n_in_8(rules_21_io_n_in_8),
    .io_n_in_9(rules_21_io_n_in_9),
    .io_n_in_10(rules_21_io_n_in_10),
    .io_n_in_11(rules_21_io_n_in_11),
    .io_n_in_12(rules_21_io_n_in_12),
    .io_n_in_13(rules_21_io_n_in_13),
    .io_n_in_14(rules_21_io_n_in_14),
    .io_n_in_15(rules_21_io_n_in_15),
    .io_n_in_16(rules_21_io_n_in_16),
    .io_n_out_0(rules_21_io_n_out_0),
    .io_n_out_1(rules_21_io_n_out_1),
    .io_n_out_2(rules_21_io_n_out_2),
    .io_n_out_3(rules_21_io_n_out_3),
    .io_n_out_4(rules_21_io_n_out_4),
    .io_n_out_5(rules_21_io_n_out_5),
    .io_n_out_6(rules_21_io_n_out_6),
    .io_n_out_7(rules_21_io_n_out_7),
    .io_n_out_8(rules_21_io_n_out_8),
    .io_n_out_9(rules_21_io_n_out_9),
    .io_n_out_10(rules_21_io_n_out_10),
    .io_n_out_11(rules_21_io_n_out_11),
    .io_n_out_12(rules_21_io_n_out_12),
    .io_n_out_13(rules_21_io_n_out_13),
    .io_n_out_14(rules_21_io_n_out_14),
    .io_n_out_15(rules_21_io_n_out_15),
    .io_n_out_16(rules_21_io_n_out_16),
    .io_x_in(rules_21_io_x_in),
    .io_x_out(rules_21_io_x_out)
  );
  Crit_5 rules_22 ( // @[system.scala 21:16]
    .io_en_r(rules_22_io_en_r),
    .io_n_in_0(rules_22_io_n_in_0),
    .io_n_in_1(rules_22_io_n_in_1),
    .io_n_in_2(rules_22_io_n_in_2),
    .io_n_in_3(rules_22_io_n_in_3),
    .io_n_in_4(rules_22_io_n_in_4),
    .io_n_in_5(rules_22_io_n_in_5),
    .io_n_in_6(rules_22_io_n_in_6),
    .io_n_in_7(rules_22_io_n_in_7),
    .io_n_in_8(rules_22_io_n_in_8),
    .io_n_in_9(rules_22_io_n_in_9),
    .io_n_in_10(rules_22_io_n_in_10),
    .io_n_in_11(rules_22_io_n_in_11),
    .io_n_in_12(rules_22_io_n_in_12),
    .io_n_in_13(rules_22_io_n_in_13),
    .io_n_in_14(rules_22_io_n_in_14),
    .io_n_in_15(rules_22_io_n_in_15),
    .io_n_in_16(rules_22_io_n_in_16),
    .io_n_out_0(rules_22_io_n_out_0),
    .io_n_out_1(rules_22_io_n_out_1),
    .io_n_out_2(rules_22_io_n_out_2),
    .io_n_out_3(rules_22_io_n_out_3),
    .io_n_out_4(rules_22_io_n_out_4),
    .io_n_out_5(rules_22_io_n_out_5),
    .io_n_out_6(rules_22_io_n_out_6),
    .io_n_out_7(rules_22_io_n_out_7),
    .io_n_out_8(rules_22_io_n_out_8),
    .io_n_out_9(rules_22_io_n_out_9),
    .io_n_out_10(rules_22_io_n_out_10),
    .io_n_out_11(rules_22_io_n_out_11),
    .io_n_out_12(rules_22_io_n_out_12),
    .io_n_out_13(rules_22_io_n_out_13),
    .io_n_out_14(rules_22_io_n_out_14),
    .io_n_out_15(rules_22_io_n_out_15),
    .io_n_out_16(rules_22_io_n_out_16),
    .io_x_in(rules_22_io_x_in),
    .io_x_out(rules_22_io_x_out)
  );
  Crit_6 rules_23 ( // @[system.scala 21:16]
    .io_en_r(rules_23_io_en_r),
    .io_n_in_0(rules_23_io_n_in_0),
    .io_n_in_1(rules_23_io_n_in_1),
    .io_n_in_2(rules_23_io_n_in_2),
    .io_n_in_3(rules_23_io_n_in_3),
    .io_n_in_4(rules_23_io_n_in_4),
    .io_n_in_5(rules_23_io_n_in_5),
    .io_n_in_6(rules_23_io_n_in_6),
    .io_n_in_7(rules_23_io_n_in_7),
    .io_n_in_8(rules_23_io_n_in_8),
    .io_n_in_9(rules_23_io_n_in_9),
    .io_n_in_10(rules_23_io_n_in_10),
    .io_n_in_11(rules_23_io_n_in_11),
    .io_n_in_12(rules_23_io_n_in_12),
    .io_n_in_13(rules_23_io_n_in_13),
    .io_n_in_14(rules_23_io_n_in_14),
    .io_n_in_15(rules_23_io_n_in_15),
    .io_n_in_16(rules_23_io_n_in_16),
    .io_n_out_0(rules_23_io_n_out_0),
    .io_n_out_1(rules_23_io_n_out_1),
    .io_n_out_2(rules_23_io_n_out_2),
    .io_n_out_3(rules_23_io_n_out_3),
    .io_n_out_4(rules_23_io_n_out_4),
    .io_n_out_5(rules_23_io_n_out_5),
    .io_n_out_6(rules_23_io_n_out_6),
    .io_n_out_7(rules_23_io_n_out_7),
    .io_n_out_8(rules_23_io_n_out_8),
    .io_n_out_9(rules_23_io_n_out_9),
    .io_n_out_10(rules_23_io_n_out_10),
    .io_n_out_11(rules_23_io_n_out_11),
    .io_n_out_12(rules_23_io_n_out_12),
    .io_n_out_13(rules_23_io_n_out_13),
    .io_n_out_14(rules_23_io_n_out_14),
    .io_n_out_15(rules_23_io_n_out_15),
    .io_n_out_16(rules_23_io_n_out_16),
    .io_x_in(rules_23_io_x_in),
    .io_x_out(rules_23_io_x_out)
  );
  Crit_7 rules_24 ( // @[system.scala 21:16]
    .io_en_r(rules_24_io_en_r),
    .io_n_in_0(rules_24_io_n_in_0),
    .io_n_in_1(rules_24_io_n_in_1),
    .io_n_in_2(rules_24_io_n_in_2),
    .io_n_in_3(rules_24_io_n_in_3),
    .io_n_in_4(rules_24_io_n_in_4),
    .io_n_in_5(rules_24_io_n_in_5),
    .io_n_in_6(rules_24_io_n_in_6),
    .io_n_in_7(rules_24_io_n_in_7),
    .io_n_in_8(rules_24_io_n_in_8),
    .io_n_in_9(rules_24_io_n_in_9),
    .io_n_in_10(rules_24_io_n_in_10),
    .io_n_in_11(rules_24_io_n_in_11),
    .io_n_in_12(rules_24_io_n_in_12),
    .io_n_in_13(rules_24_io_n_in_13),
    .io_n_in_14(rules_24_io_n_in_14),
    .io_n_in_15(rules_24_io_n_in_15),
    .io_n_in_16(rules_24_io_n_in_16),
    .io_n_out_0(rules_24_io_n_out_0),
    .io_n_out_1(rules_24_io_n_out_1),
    .io_n_out_2(rules_24_io_n_out_2),
    .io_n_out_3(rules_24_io_n_out_3),
    .io_n_out_4(rules_24_io_n_out_4),
    .io_n_out_5(rules_24_io_n_out_5),
    .io_n_out_6(rules_24_io_n_out_6),
    .io_n_out_7(rules_24_io_n_out_7),
    .io_n_out_8(rules_24_io_n_out_8),
    .io_n_out_9(rules_24_io_n_out_9),
    .io_n_out_10(rules_24_io_n_out_10),
    .io_n_out_11(rules_24_io_n_out_11),
    .io_n_out_12(rules_24_io_n_out_12),
    .io_n_out_13(rules_24_io_n_out_13),
    .io_n_out_14(rules_24_io_n_out_14),
    .io_n_out_15(rules_24_io_n_out_15),
    .io_n_out_16(rules_24_io_n_out_16),
    .io_x_in(rules_24_io_x_in),
    .io_x_out(rules_24_io_x_out)
  );
  Crit_8 rules_25 ( // @[system.scala 21:16]
    .io_en_r(rules_25_io_en_r),
    .io_n_in_0(rules_25_io_n_in_0),
    .io_n_in_1(rules_25_io_n_in_1),
    .io_n_in_2(rules_25_io_n_in_2),
    .io_n_in_3(rules_25_io_n_in_3),
    .io_n_in_4(rules_25_io_n_in_4),
    .io_n_in_5(rules_25_io_n_in_5),
    .io_n_in_6(rules_25_io_n_in_6),
    .io_n_in_7(rules_25_io_n_in_7),
    .io_n_in_8(rules_25_io_n_in_8),
    .io_n_in_9(rules_25_io_n_in_9),
    .io_n_in_10(rules_25_io_n_in_10),
    .io_n_in_11(rules_25_io_n_in_11),
    .io_n_in_12(rules_25_io_n_in_12),
    .io_n_in_13(rules_25_io_n_in_13),
    .io_n_in_14(rules_25_io_n_in_14),
    .io_n_in_15(rules_25_io_n_in_15),
    .io_n_in_16(rules_25_io_n_in_16),
    .io_n_out_0(rules_25_io_n_out_0),
    .io_n_out_1(rules_25_io_n_out_1),
    .io_n_out_2(rules_25_io_n_out_2),
    .io_n_out_3(rules_25_io_n_out_3),
    .io_n_out_4(rules_25_io_n_out_4),
    .io_n_out_5(rules_25_io_n_out_5),
    .io_n_out_6(rules_25_io_n_out_6),
    .io_n_out_7(rules_25_io_n_out_7),
    .io_n_out_8(rules_25_io_n_out_8),
    .io_n_out_9(rules_25_io_n_out_9),
    .io_n_out_10(rules_25_io_n_out_10),
    .io_n_out_11(rules_25_io_n_out_11),
    .io_n_out_12(rules_25_io_n_out_12),
    .io_n_out_13(rules_25_io_n_out_13),
    .io_n_out_14(rules_25_io_n_out_14),
    .io_n_out_15(rules_25_io_n_out_15),
    .io_n_out_16(rules_25_io_n_out_16),
    .io_x_in(rules_25_io_x_in),
    .io_x_out(rules_25_io_x_out)
  );
  Crit_9 rules_26 ( // @[system.scala 21:16]
    .io_en_r(rules_26_io_en_r),
    .io_n_in_0(rules_26_io_n_in_0),
    .io_n_in_1(rules_26_io_n_in_1),
    .io_n_in_2(rules_26_io_n_in_2),
    .io_n_in_3(rules_26_io_n_in_3),
    .io_n_in_4(rules_26_io_n_in_4),
    .io_n_in_5(rules_26_io_n_in_5),
    .io_n_in_6(rules_26_io_n_in_6),
    .io_n_in_7(rules_26_io_n_in_7),
    .io_n_in_8(rules_26_io_n_in_8),
    .io_n_in_9(rules_26_io_n_in_9),
    .io_n_in_10(rules_26_io_n_in_10),
    .io_n_in_11(rules_26_io_n_in_11),
    .io_n_in_12(rules_26_io_n_in_12),
    .io_n_in_13(rules_26_io_n_in_13),
    .io_n_in_14(rules_26_io_n_in_14),
    .io_n_in_15(rules_26_io_n_in_15),
    .io_n_in_16(rules_26_io_n_in_16),
    .io_n_out_0(rules_26_io_n_out_0),
    .io_n_out_1(rules_26_io_n_out_1),
    .io_n_out_2(rules_26_io_n_out_2),
    .io_n_out_3(rules_26_io_n_out_3),
    .io_n_out_4(rules_26_io_n_out_4),
    .io_n_out_5(rules_26_io_n_out_5),
    .io_n_out_6(rules_26_io_n_out_6),
    .io_n_out_7(rules_26_io_n_out_7),
    .io_n_out_8(rules_26_io_n_out_8),
    .io_n_out_9(rules_26_io_n_out_9),
    .io_n_out_10(rules_26_io_n_out_10),
    .io_n_out_11(rules_26_io_n_out_11),
    .io_n_out_12(rules_26_io_n_out_12),
    .io_n_out_13(rules_26_io_n_out_13),
    .io_n_out_14(rules_26_io_n_out_14),
    .io_n_out_15(rules_26_io_n_out_15),
    .io_n_out_16(rules_26_io_n_out_16),
    .io_x_in(rules_26_io_x_in),
    .io_x_out(rules_26_io_x_out)
  );
  Crit_10 rules_27 ( // @[system.scala 21:16]
    .io_en_r(rules_27_io_en_r),
    .io_n_in_0(rules_27_io_n_in_0),
    .io_n_in_1(rules_27_io_n_in_1),
    .io_n_in_2(rules_27_io_n_in_2),
    .io_n_in_3(rules_27_io_n_in_3),
    .io_n_in_4(rules_27_io_n_in_4),
    .io_n_in_5(rules_27_io_n_in_5),
    .io_n_in_6(rules_27_io_n_in_6),
    .io_n_in_7(rules_27_io_n_in_7),
    .io_n_in_8(rules_27_io_n_in_8),
    .io_n_in_9(rules_27_io_n_in_9),
    .io_n_in_10(rules_27_io_n_in_10),
    .io_n_in_11(rules_27_io_n_in_11),
    .io_n_in_12(rules_27_io_n_in_12),
    .io_n_in_13(rules_27_io_n_in_13),
    .io_n_in_14(rules_27_io_n_in_14),
    .io_n_in_15(rules_27_io_n_in_15),
    .io_n_in_16(rules_27_io_n_in_16),
    .io_n_out_0(rules_27_io_n_out_0),
    .io_n_out_1(rules_27_io_n_out_1),
    .io_n_out_2(rules_27_io_n_out_2),
    .io_n_out_3(rules_27_io_n_out_3),
    .io_n_out_4(rules_27_io_n_out_4),
    .io_n_out_5(rules_27_io_n_out_5),
    .io_n_out_6(rules_27_io_n_out_6),
    .io_n_out_7(rules_27_io_n_out_7),
    .io_n_out_8(rules_27_io_n_out_8),
    .io_n_out_9(rules_27_io_n_out_9),
    .io_n_out_10(rules_27_io_n_out_10),
    .io_n_out_11(rules_27_io_n_out_11),
    .io_n_out_12(rules_27_io_n_out_12),
    .io_n_out_13(rules_27_io_n_out_13),
    .io_n_out_14(rules_27_io_n_out_14),
    .io_n_out_15(rules_27_io_n_out_15),
    .io_n_out_16(rules_27_io_n_out_16),
    .io_x_in(rules_27_io_x_in),
    .io_x_out(rules_27_io_x_out)
  );
  Crit_11 rules_28 ( // @[system.scala 21:16]
    .io_en_r(rules_28_io_en_r),
    .io_n_in_0(rules_28_io_n_in_0),
    .io_n_in_1(rules_28_io_n_in_1),
    .io_n_in_2(rules_28_io_n_in_2),
    .io_n_in_3(rules_28_io_n_in_3),
    .io_n_in_4(rules_28_io_n_in_4),
    .io_n_in_5(rules_28_io_n_in_5),
    .io_n_in_6(rules_28_io_n_in_6),
    .io_n_in_7(rules_28_io_n_in_7),
    .io_n_in_8(rules_28_io_n_in_8),
    .io_n_in_9(rules_28_io_n_in_9),
    .io_n_in_10(rules_28_io_n_in_10),
    .io_n_in_11(rules_28_io_n_in_11),
    .io_n_in_12(rules_28_io_n_in_12),
    .io_n_in_13(rules_28_io_n_in_13),
    .io_n_in_14(rules_28_io_n_in_14),
    .io_n_in_15(rules_28_io_n_in_15),
    .io_n_in_16(rules_28_io_n_in_16),
    .io_n_out_0(rules_28_io_n_out_0),
    .io_n_out_1(rules_28_io_n_out_1),
    .io_n_out_2(rules_28_io_n_out_2),
    .io_n_out_3(rules_28_io_n_out_3),
    .io_n_out_4(rules_28_io_n_out_4),
    .io_n_out_5(rules_28_io_n_out_5),
    .io_n_out_6(rules_28_io_n_out_6),
    .io_n_out_7(rules_28_io_n_out_7),
    .io_n_out_8(rules_28_io_n_out_8),
    .io_n_out_9(rules_28_io_n_out_9),
    .io_n_out_10(rules_28_io_n_out_10),
    .io_n_out_11(rules_28_io_n_out_11),
    .io_n_out_12(rules_28_io_n_out_12),
    .io_n_out_13(rules_28_io_n_out_13),
    .io_n_out_14(rules_28_io_n_out_14),
    .io_n_out_15(rules_28_io_n_out_15),
    .io_n_out_16(rules_28_io_n_out_16),
    .io_x_in(rules_28_io_x_in),
    .io_x_out(rules_28_io_x_out)
  );
  Crit_12 rules_29 ( // @[system.scala 21:16]
    .io_en_r(rules_29_io_en_r),
    .io_n_in_0(rules_29_io_n_in_0),
    .io_n_in_1(rules_29_io_n_in_1),
    .io_n_in_2(rules_29_io_n_in_2),
    .io_n_in_3(rules_29_io_n_in_3),
    .io_n_in_4(rules_29_io_n_in_4),
    .io_n_in_5(rules_29_io_n_in_5),
    .io_n_in_6(rules_29_io_n_in_6),
    .io_n_in_7(rules_29_io_n_in_7),
    .io_n_in_8(rules_29_io_n_in_8),
    .io_n_in_9(rules_29_io_n_in_9),
    .io_n_in_10(rules_29_io_n_in_10),
    .io_n_in_11(rules_29_io_n_in_11),
    .io_n_in_12(rules_29_io_n_in_12),
    .io_n_in_13(rules_29_io_n_in_13),
    .io_n_in_14(rules_29_io_n_in_14),
    .io_n_in_15(rules_29_io_n_in_15),
    .io_n_in_16(rules_29_io_n_in_16),
    .io_n_out_0(rules_29_io_n_out_0),
    .io_n_out_1(rules_29_io_n_out_1),
    .io_n_out_2(rules_29_io_n_out_2),
    .io_n_out_3(rules_29_io_n_out_3),
    .io_n_out_4(rules_29_io_n_out_4),
    .io_n_out_5(rules_29_io_n_out_5),
    .io_n_out_6(rules_29_io_n_out_6),
    .io_n_out_7(rules_29_io_n_out_7),
    .io_n_out_8(rules_29_io_n_out_8),
    .io_n_out_9(rules_29_io_n_out_9),
    .io_n_out_10(rules_29_io_n_out_10),
    .io_n_out_11(rules_29_io_n_out_11),
    .io_n_out_12(rules_29_io_n_out_12),
    .io_n_out_13(rules_29_io_n_out_13),
    .io_n_out_14(rules_29_io_n_out_14),
    .io_n_out_15(rules_29_io_n_out_15),
    .io_n_out_16(rules_29_io_n_out_16),
    .io_x_in(rules_29_io_x_in),
    .io_x_out(rules_29_io_x_out)
  );
  Crit_13 rules_30 ( // @[system.scala 21:16]
    .io_en_r(rules_30_io_en_r),
    .io_n_in_0(rules_30_io_n_in_0),
    .io_n_in_1(rules_30_io_n_in_1),
    .io_n_in_2(rules_30_io_n_in_2),
    .io_n_in_3(rules_30_io_n_in_3),
    .io_n_in_4(rules_30_io_n_in_4),
    .io_n_in_5(rules_30_io_n_in_5),
    .io_n_in_6(rules_30_io_n_in_6),
    .io_n_in_7(rules_30_io_n_in_7),
    .io_n_in_8(rules_30_io_n_in_8),
    .io_n_in_9(rules_30_io_n_in_9),
    .io_n_in_10(rules_30_io_n_in_10),
    .io_n_in_11(rules_30_io_n_in_11),
    .io_n_in_12(rules_30_io_n_in_12),
    .io_n_in_13(rules_30_io_n_in_13),
    .io_n_in_14(rules_30_io_n_in_14),
    .io_n_in_15(rules_30_io_n_in_15),
    .io_n_in_16(rules_30_io_n_in_16),
    .io_n_out_0(rules_30_io_n_out_0),
    .io_n_out_1(rules_30_io_n_out_1),
    .io_n_out_2(rules_30_io_n_out_2),
    .io_n_out_3(rules_30_io_n_out_3),
    .io_n_out_4(rules_30_io_n_out_4),
    .io_n_out_5(rules_30_io_n_out_5),
    .io_n_out_6(rules_30_io_n_out_6),
    .io_n_out_7(rules_30_io_n_out_7),
    .io_n_out_8(rules_30_io_n_out_8),
    .io_n_out_9(rules_30_io_n_out_9),
    .io_n_out_10(rules_30_io_n_out_10),
    .io_n_out_11(rules_30_io_n_out_11),
    .io_n_out_12(rules_30_io_n_out_12),
    .io_n_out_13(rules_30_io_n_out_13),
    .io_n_out_14(rules_30_io_n_out_14),
    .io_n_out_15(rules_30_io_n_out_15),
    .io_n_out_16(rules_30_io_n_out_16),
    .io_x_in(rules_30_io_x_in),
    .io_x_out(rules_30_io_x_out)
  );
  Crit_14 rules_31 ( // @[system.scala 21:16]
    .io_en_r(rules_31_io_en_r),
    .io_n_in_0(rules_31_io_n_in_0),
    .io_n_in_1(rules_31_io_n_in_1),
    .io_n_in_2(rules_31_io_n_in_2),
    .io_n_in_3(rules_31_io_n_in_3),
    .io_n_in_4(rules_31_io_n_in_4),
    .io_n_in_5(rules_31_io_n_in_5),
    .io_n_in_6(rules_31_io_n_in_6),
    .io_n_in_7(rules_31_io_n_in_7),
    .io_n_in_8(rules_31_io_n_in_8),
    .io_n_in_9(rules_31_io_n_in_9),
    .io_n_in_10(rules_31_io_n_in_10),
    .io_n_in_11(rules_31_io_n_in_11),
    .io_n_in_12(rules_31_io_n_in_12),
    .io_n_in_13(rules_31_io_n_in_13),
    .io_n_in_14(rules_31_io_n_in_14),
    .io_n_in_15(rules_31_io_n_in_15),
    .io_n_in_16(rules_31_io_n_in_16),
    .io_n_out_0(rules_31_io_n_out_0),
    .io_n_out_1(rules_31_io_n_out_1),
    .io_n_out_2(rules_31_io_n_out_2),
    .io_n_out_3(rules_31_io_n_out_3),
    .io_n_out_4(rules_31_io_n_out_4),
    .io_n_out_5(rules_31_io_n_out_5),
    .io_n_out_6(rules_31_io_n_out_6),
    .io_n_out_7(rules_31_io_n_out_7),
    .io_n_out_8(rules_31_io_n_out_8),
    .io_n_out_9(rules_31_io_n_out_9),
    .io_n_out_10(rules_31_io_n_out_10),
    .io_n_out_11(rules_31_io_n_out_11),
    .io_n_out_12(rules_31_io_n_out_12),
    .io_n_out_13(rules_31_io_n_out_13),
    .io_n_out_14(rules_31_io_n_out_14),
    .io_n_out_15(rules_31_io_n_out_15),
    .io_n_out_16(rules_31_io_n_out_16),
    .io_x_in(rules_31_io_x_in),
    .io_x_out(rules_31_io_x_out)
  );
  Crit_15 rules_32 ( // @[system.scala 21:16]
    .io_en_r(rules_32_io_en_r),
    .io_n_in_0(rules_32_io_n_in_0),
    .io_n_in_1(rules_32_io_n_in_1),
    .io_n_in_2(rules_32_io_n_in_2),
    .io_n_in_3(rules_32_io_n_in_3),
    .io_n_in_4(rules_32_io_n_in_4),
    .io_n_in_5(rules_32_io_n_in_5),
    .io_n_in_6(rules_32_io_n_in_6),
    .io_n_in_7(rules_32_io_n_in_7),
    .io_n_in_8(rules_32_io_n_in_8),
    .io_n_in_9(rules_32_io_n_in_9),
    .io_n_in_10(rules_32_io_n_in_10),
    .io_n_in_11(rules_32_io_n_in_11),
    .io_n_in_12(rules_32_io_n_in_12),
    .io_n_in_13(rules_32_io_n_in_13),
    .io_n_in_14(rules_32_io_n_in_14),
    .io_n_in_15(rules_32_io_n_in_15),
    .io_n_in_16(rules_32_io_n_in_16),
    .io_n_out_0(rules_32_io_n_out_0),
    .io_n_out_1(rules_32_io_n_out_1),
    .io_n_out_2(rules_32_io_n_out_2),
    .io_n_out_3(rules_32_io_n_out_3),
    .io_n_out_4(rules_32_io_n_out_4),
    .io_n_out_5(rules_32_io_n_out_5),
    .io_n_out_6(rules_32_io_n_out_6),
    .io_n_out_7(rules_32_io_n_out_7),
    .io_n_out_8(rules_32_io_n_out_8),
    .io_n_out_9(rules_32_io_n_out_9),
    .io_n_out_10(rules_32_io_n_out_10),
    .io_n_out_11(rules_32_io_n_out_11),
    .io_n_out_12(rules_32_io_n_out_12),
    .io_n_out_13(rules_32_io_n_out_13),
    .io_n_out_14(rules_32_io_n_out_14),
    .io_n_out_15(rules_32_io_n_out_15),
    .io_n_out_16(rules_32_io_n_out_16),
    .io_x_in(rules_32_io_x_in),
    .io_x_out(rules_32_io_x_out)
  );
  Exit rules_33 ( // @[system.scala 24:16]
    .io_en_r(rules_33_io_en_r),
    .io_n_in_0(rules_33_io_n_in_0),
    .io_n_in_1(rules_33_io_n_in_1),
    .io_n_in_2(rules_33_io_n_in_2),
    .io_n_in_3(rules_33_io_n_in_3),
    .io_n_in_4(rules_33_io_n_in_4),
    .io_n_in_5(rules_33_io_n_in_5),
    .io_n_in_6(rules_33_io_n_in_6),
    .io_n_in_7(rules_33_io_n_in_7),
    .io_n_in_8(rules_33_io_n_in_8),
    .io_n_in_9(rules_33_io_n_in_9),
    .io_n_in_10(rules_33_io_n_in_10),
    .io_n_in_11(rules_33_io_n_in_11),
    .io_n_in_12(rules_33_io_n_in_12),
    .io_n_in_13(rules_33_io_n_in_13),
    .io_n_in_14(rules_33_io_n_in_14),
    .io_n_in_15(rules_33_io_n_in_15),
    .io_n_in_16(rules_33_io_n_in_16),
    .io_n_out_0(rules_33_io_n_out_0),
    .io_n_out_1(rules_33_io_n_out_1),
    .io_n_out_2(rules_33_io_n_out_2),
    .io_n_out_3(rules_33_io_n_out_3),
    .io_n_out_4(rules_33_io_n_out_4),
    .io_n_out_5(rules_33_io_n_out_5),
    .io_n_out_6(rules_33_io_n_out_6),
    .io_n_out_7(rules_33_io_n_out_7),
    .io_n_out_8(rules_33_io_n_out_8),
    .io_n_out_9(rules_33_io_n_out_9),
    .io_n_out_10(rules_33_io_n_out_10),
    .io_n_out_11(rules_33_io_n_out_11),
    .io_n_out_12(rules_33_io_n_out_12),
    .io_n_out_13(rules_33_io_n_out_13),
    .io_n_out_14(rules_33_io_n_out_14),
    .io_n_out_15(rules_33_io_n_out_15),
    .io_n_out_16(rules_33_io_n_out_16),
    .io_x_in(rules_33_io_x_in),
    .io_x_out(rules_33_io_x_out)
  );
  Exit_1 rules_34 ( // @[system.scala 24:16]
    .io_en_r(rules_34_io_en_r),
    .io_n_in_0(rules_34_io_n_in_0),
    .io_n_in_1(rules_34_io_n_in_1),
    .io_n_in_2(rules_34_io_n_in_2),
    .io_n_in_3(rules_34_io_n_in_3),
    .io_n_in_4(rules_34_io_n_in_4),
    .io_n_in_5(rules_34_io_n_in_5),
    .io_n_in_6(rules_34_io_n_in_6),
    .io_n_in_7(rules_34_io_n_in_7),
    .io_n_in_8(rules_34_io_n_in_8),
    .io_n_in_9(rules_34_io_n_in_9),
    .io_n_in_10(rules_34_io_n_in_10),
    .io_n_in_11(rules_34_io_n_in_11),
    .io_n_in_12(rules_34_io_n_in_12),
    .io_n_in_13(rules_34_io_n_in_13),
    .io_n_in_14(rules_34_io_n_in_14),
    .io_n_in_15(rules_34_io_n_in_15),
    .io_n_in_16(rules_34_io_n_in_16),
    .io_n_out_0(rules_34_io_n_out_0),
    .io_n_out_1(rules_34_io_n_out_1),
    .io_n_out_2(rules_34_io_n_out_2),
    .io_n_out_3(rules_34_io_n_out_3),
    .io_n_out_4(rules_34_io_n_out_4),
    .io_n_out_5(rules_34_io_n_out_5),
    .io_n_out_6(rules_34_io_n_out_6),
    .io_n_out_7(rules_34_io_n_out_7),
    .io_n_out_8(rules_34_io_n_out_8),
    .io_n_out_9(rules_34_io_n_out_9),
    .io_n_out_10(rules_34_io_n_out_10),
    .io_n_out_11(rules_34_io_n_out_11),
    .io_n_out_12(rules_34_io_n_out_12),
    .io_n_out_13(rules_34_io_n_out_13),
    .io_n_out_14(rules_34_io_n_out_14),
    .io_n_out_15(rules_34_io_n_out_15),
    .io_n_out_16(rules_34_io_n_out_16),
    .io_x_in(rules_34_io_x_in),
    .io_x_out(rules_34_io_x_out)
  );
  Exit_2 rules_35 ( // @[system.scala 24:16]
    .io_en_r(rules_35_io_en_r),
    .io_n_in_0(rules_35_io_n_in_0),
    .io_n_in_1(rules_35_io_n_in_1),
    .io_n_in_2(rules_35_io_n_in_2),
    .io_n_in_3(rules_35_io_n_in_3),
    .io_n_in_4(rules_35_io_n_in_4),
    .io_n_in_5(rules_35_io_n_in_5),
    .io_n_in_6(rules_35_io_n_in_6),
    .io_n_in_7(rules_35_io_n_in_7),
    .io_n_in_8(rules_35_io_n_in_8),
    .io_n_in_9(rules_35_io_n_in_9),
    .io_n_in_10(rules_35_io_n_in_10),
    .io_n_in_11(rules_35_io_n_in_11),
    .io_n_in_12(rules_35_io_n_in_12),
    .io_n_in_13(rules_35_io_n_in_13),
    .io_n_in_14(rules_35_io_n_in_14),
    .io_n_in_15(rules_35_io_n_in_15),
    .io_n_in_16(rules_35_io_n_in_16),
    .io_n_out_0(rules_35_io_n_out_0),
    .io_n_out_1(rules_35_io_n_out_1),
    .io_n_out_2(rules_35_io_n_out_2),
    .io_n_out_3(rules_35_io_n_out_3),
    .io_n_out_4(rules_35_io_n_out_4),
    .io_n_out_5(rules_35_io_n_out_5),
    .io_n_out_6(rules_35_io_n_out_6),
    .io_n_out_7(rules_35_io_n_out_7),
    .io_n_out_8(rules_35_io_n_out_8),
    .io_n_out_9(rules_35_io_n_out_9),
    .io_n_out_10(rules_35_io_n_out_10),
    .io_n_out_11(rules_35_io_n_out_11),
    .io_n_out_12(rules_35_io_n_out_12),
    .io_n_out_13(rules_35_io_n_out_13),
    .io_n_out_14(rules_35_io_n_out_14),
    .io_n_out_15(rules_35_io_n_out_15),
    .io_n_out_16(rules_35_io_n_out_16),
    .io_x_in(rules_35_io_x_in),
    .io_x_out(rules_35_io_x_out)
  );
  Exit_3 rules_36 ( // @[system.scala 24:16]
    .io_en_r(rules_36_io_en_r),
    .io_n_in_0(rules_36_io_n_in_0),
    .io_n_in_1(rules_36_io_n_in_1),
    .io_n_in_2(rules_36_io_n_in_2),
    .io_n_in_3(rules_36_io_n_in_3),
    .io_n_in_4(rules_36_io_n_in_4),
    .io_n_in_5(rules_36_io_n_in_5),
    .io_n_in_6(rules_36_io_n_in_6),
    .io_n_in_7(rules_36_io_n_in_7),
    .io_n_in_8(rules_36_io_n_in_8),
    .io_n_in_9(rules_36_io_n_in_9),
    .io_n_in_10(rules_36_io_n_in_10),
    .io_n_in_11(rules_36_io_n_in_11),
    .io_n_in_12(rules_36_io_n_in_12),
    .io_n_in_13(rules_36_io_n_in_13),
    .io_n_in_14(rules_36_io_n_in_14),
    .io_n_in_15(rules_36_io_n_in_15),
    .io_n_in_16(rules_36_io_n_in_16),
    .io_n_out_0(rules_36_io_n_out_0),
    .io_n_out_1(rules_36_io_n_out_1),
    .io_n_out_2(rules_36_io_n_out_2),
    .io_n_out_3(rules_36_io_n_out_3),
    .io_n_out_4(rules_36_io_n_out_4),
    .io_n_out_5(rules_36_io_n_out_5),
    .io_n_out_6(rules_36_io_n_out_6),
    .io_n_out_7(rules_36_io_n_out_7),
    .io_n_out_8(rules_36_io_n_out_8),
    .io_n_out_9(rules_36_io_n_out_9),
    .io_n_out_10(rules_36_io_n_out_10),
    .io_n_out_11(rules_36_io_n_out_11),
    .io_n_out_12(rules_36_io_n_out_12),
    .io_n_out_13(rules_36_io_n_out_13),
    .io_n_out_14(rules_36_io_n_out_14),
    .io_n_out_15(rules_36_io_n_out_15),
    .io_n_out_16(rules_36_io_n_out_16),
    .io_x_in(rules_36_io_x_in),
    .io_x_out(rules_36_io_x_out)
  );
  Exit_4 rules_37 ( // @[system.scala 24:16]
    .io_en_r(rules_37_io_en_r),
    .io_n_in_0(rules_37_io_n_in_0),
    .io_n_in_1(rules_37_io_n_in_1),
    .io_n_in_2(rules_37_io_n_in_2),
    .io_n_in_3(rules_37_io_n_in_3),
    .io_n_in_4(rules_37_io_n_in_4),
    .io_n_in_5(rules_37_io_n_in_5),
    .io_n_in_6(rules_37_io_n_in_6),
    .io_n_in_7(rules_37_io_n_in_7),
    .io_n_in_8(rules_37_io_n_in_8),
    .io_n_in_9(rules_37_io_n_in_9),
    .io_n_in_10(rules_37_io_n_in_10),
    .io_n_in_11(rules_37_io_n_in_11),
    .io_n_in_12(rules_37_io_n_in_12),
    .io_n_in_13(rules_37_io_n_in_13),
    .io_n_in_14(rules_37_io_n_in_14),
    .io_n_in_15(rules_37_io_n_in_15),
    .io_n_in_16(rules_37_io_n_in_16),
    .io_n_out_0(rules_37_io_n_out_0),
    .io_n_out_1(rules_37_io_n_out_1),
    .io_n_out_2(rules_37_io_n_out_2),
    .io_n_out_3(rules_37_io_n_out_3),
    .io_n_out_4(rules_37_io_n_out_4),
    .io_n_out_5(rules_37_io_n_out_5),
    .io_n_out_6(rules_37_io_n_out_6),
    .io_n_out_7(rules_37_io_n_out_7),
    .io_n_out_8(rules_37_io_n_out_8),
    .io_n_out_9(rules_37_io_n_out_9),
    .io_n_out_10(rules_37_io_n_out_10),
    .io_n_out_11(rules_37_io_n_out_11),
    .io_n_out_12(rules_37_io_n_out_12),
    .io_n_out_13(rules_37_io_n_out_13),
    .io_n_out_14(rules_37_io_n_out_14),
    .io_n_out_15(rules_37_io_n_out_15),
    .io_n_out_16(rules_37_io_n_out_16),
    .io_x_in(rules_37_io_x_in),
    .io_x_out(rules_37_io_x_out)
  );
  Exit_5 rules_38 ( // @[system.scala 24:16]
    .io_en_r(rules_38_io_en_r),
    .io_n_in_0(rules_38_io_n_in_0),
    .io_n_in_1(rules_38_io_n_in_1),
    .io_n_in_2(rules_38_io_n_in_2),
    .io_n_in_3(rules_38_io_n_in_3),
    .io_n_in_4(rules_38_io_n_in_4),
    .io_n_in_5(rules_38_io_n_in_5),
    .io_n_in_6(rules_38_io_n_in_6),
    .io_n_in_7(rules_38_io_n_in_7),
    .io_n_in_8(rules_38_io_n_in_8),
    .io_n_in_9(rules_38_io_n_in_9),
    .io_n_in_10(rules_38_io_n_in_10),
    .io_n_in_11(rules_38_io_n_in_11),
    .io_n_in_12(rules_38_io_n_in_12),
    .io_n_in_13(rules_38_io_n_in_13),
    .io_n_in_14(rules_38_io_n_in_14),
    .io_n_in_15(rules_38_io_n_in_15),
    .io_n_in_16(rules_38_io_n_in_16),
    .io_n_out_0(rules_38_io_n_out_0),
    .io_n_out_1(rules_38_io_n_out_1),
    .io_n_out_2(rules_38_io_n_out_2),
    .io_n_out_3(rules_38_io_n_out_3),
    .io_n_out_4(rules_38_io_n_out_4),
    .io_n_out_5(rules_38_io_n_out_5),
    .io_n_out_6(rules_38_io_n_out_6),
    .io_n_out_7(rules_38_io_n_out_7),
    .io_n_out_8(rules_38_io_n_out_8),
    .io_n_out_9(rules_38_io_n_out_9),
    .io_n_out_10(rules_38_io_n_out_10),
    .io_n_out_11(rules_38_io_n_out_11),
    .io_n_out_12(rules_38_io_n_out_12),
    .io_n_out_13(rules_38_io_n_out_13),
    .io_n_out_14(rules_38_io_n_out_14),
    .io_n_out_15(rules_38_io_n_out_15),
    .io_n_out_16(rules_38_io_n_out_16),
    .io_x_in(rules_38_io_x_in),
    .io_x_out(rules_38_io_x_out)
  );
  Exit_6 rules_39 ( // @[system.scala 24:16]
    .io_en_r(rules_39_io_en_r),
    .io_n_in_0(rules_39_io_n_in_0),
    .io_n_in_1(rules_39_io_n_in_1),
    .io_n_in_2(rules_39_io_n_in_2),
    .io_n_in_3(rules_39_io_n_in_3),
    .io_n_in_4(rules_39_io_n_in_4),
    .io_n_in_5(rules_39_io_n_in_5),
    .io_n_in_6(rules_39_io_n_in_6),
    .io_n_in_7(rules_39_io_n_in_7),
    .io_n_in_8(rules_39_io_n_in_8),
    .io_n_in_9(rules_39_io_n_in_9),
    .io_n_in_10(rules_39_io_n_in_10),
    .io_n_in_11(rules_39_io_n_in_11),
    .io_n_in_12(rules_39_io_n_in_12),
    .io_n_in_13(rules_39_io_n_in_13),
    .io_n_in_14(rules_39_io_n_in_14),
    .io_n_in_15(rules_39_io_n_in_15),
    .io_n_in_16(rules_39_io_n_in_16),
    .io_n_out_0(rules_39_io_n_out_0),
    .io_n_out_1(rules_39_io_n_out_1),
    .io_n_out_2(rules_39_io_n_out_2),
    .io_n_out_3(rules_39_io_n_out_3),
    .io_n_out_4(rules_39_io_n_out_4),
    .io_n_out_5(rules_39_io_n_out_5),
    .io_n_out_6(rules_39_io_n_out_6),
    .io_n_out_7(rules_39_io_n_out_7),
    .io_n_out_8(rules_39_io_n_out_8),
    .io_n_out_9(rules_39_io_n_out_9),
    .io_n_out_10(rules_39_io_n_out_10),
    .io_n_out_11(rules_39_io_n_out_11),
    .io_n_out_12(rules_39_io_n_out_12),
    .io_n_out_13(rules_39_io_n_out_13),
    .io_n_out_14(rules_39_io_n_out_14),
    .io_n_out_15(rules_39_io_n_out_15),
    .io_n_out_16(rules_39_io_n_out_16),
    .io_x_in(rules_39_io_x_in),
    .io_x_out(rules_39_io_x_out)
  );
  Exit_7 rules_40 ( // @[system.scala 24:16]
    .io_en_r(rules_40_io_en_r),
    .io_n_in_0(rules_40_io_n_in_0),
    .io_n_in_1(rules_40_io_n_in_1),
    .io_n_in_2(rules_40_io_n_in_2),
    .io_n_in_3(rules_40_io_n_in_3),
    .io_n_in_4(rules_40_io_n_in_4),
    .io_n_in_5(rules_40_io_n_in_5),
    .io_n_in_6(rules_40_io_n_in_6),
    .io_n_in_7(rules_40_io_n_in_7),
    .io_n_in_8(rules_40_io_n_in_8),
    .io_n_in_9(rules_40_io_n_in_9),
    .io_n_in_10(rules_40_io_n_in_10),
    .io_n_in_11(rules_40_io_n_in_11),
    .io_n_in_12(rules_40_io_n_in_12),
    .io_n_in_13(rules_40_io_n_in_13),
    .io_n_in_14(rules_40_io_n_in_14),
    .io_n_in_15(rules_40_io_n_in_15),
    .io_n_in_16(rules_40_io_n_in_16),
    .io_n_out_0(rules_40_io_n_out_0),
    .io_n_out_1(rules_40_io_n_out_1),
    .io_n_out_2(rules_40_io_n_out_2),
    .io_n_out_3(rules_40_io_n_out_3),
    .io_n_out_4(rules_40_io_n_out_4),
    .io_n_out_5(rules_40_io_n_out_5),
    .io_n_out_6(rules_40_io_n_out_6),
    .io_n_out_7(rules_40_io_n_out_7),
    .io_n_out_8(rules_40_io_n_out_8),
    .io_n_out_9(rules_40_io_n_out_9),
    .io_n_out_10(rules_40_io_n_out_10),
    .io_n_out_11(rules_40_io_n_out_11),
    .io_n_out_12(rules_40_io_n_out_12),
    .io_n_out_13(rules_40_io_n_out_13),
    .io_n_out_14(rules_40_io_n_out_14),
    .io_n_out_15(rules_40_io_n_out_15),
    .io_n_out_16(rules_40_io_n_out_16),
    .io_x_in(rules_40_io_x_in),
    .io_x_out(rules_40_io_x_out)
  );
  Exit_8 rules_41 ( // @[system.scala 24:16]
    .io_en_r(rules_41_io_en_r),
    .io_n_in_0(rules_41_io_n_in_0),
    .io_n_in_1(rules_41_io_n_in_1),
    .io_n_in_2(rules_41_io_n_in_2),
    .io_n_in_3(rules_41_io_n_in_3),
    .io_n_in_4(rules_41_io_n_in_4),
    .io_n_in_5(rules_41_io_n_in_5),
    .io_n_in_6(rules_41_io_n_in_6),
    .io_n_in_7(rules_41_io_n_in_7),
    .io_n_in_8(rules_41_io_n_in_8),
    .io_n_in_9(rules_41_io_n_in_9),
    .io_n_in_10(rules_41_io_n_in_10),
    .io_n_in_11(rules_41_io_n_in_11),
    .io_n_in_12(rules_41_io_n_in_12),
    .io_n_in_13(rules_41_io_n_in_13),
    .io_n_in_14(rules_41_io_n_in_14),
    .io_n_in_15(rules_41_io_n_in_15),
    .io_n_in_16(rules_41_io_n_in_16),
    .io_n_out_0(rules_41_io_n_out_0),
    .io_n_out_1(rules_41_io_n_out_1),
    .io_n_out_2(rules_41_io_n_out_2),
    .io_n_out_3(rules_41_io_n_out_3),
    .io_n_out_4(rules_41_io_n_out_4),
    .io_n_out_5(rules_41_io_n_out_5),
    .io_n_out_6(rules_41_io_n_out_6),
    .io_n_out_7(rules_41_io_n_out_7),
    .io_n_out_8(rules_41_io_n_out_8),
    .io_n_out_9(rules_41_io_n_out_9),
    .io_n_out_10(rules_41_io_n_out_10),
    .io_n_out_11(rules_41_io_n_out_11),
    .io_n_out_12(rules_41_io_n_out_12),
    .io_n_out_13(rules_41_io_n_out_13),
    .io_n_out_14(rules_41_io_n_out_14),
    .io_n_out_15(rules_41_io_n_out_15),
    .io_n_out_16(rules_41_io_n_out_16),
    .io_x_in(rules_41_io_x_in),
    .io_x_out(rules_41_io_x_out)
  );
  Exit_9 rules_42 ( // @[system.scala 24:16]
    .io_en_r(rules_42_io_en_r),
    .io_n_in_0(rules_42_io_n_in_0),
    .io_n_in_1(rules_42_io_n_in_1),
    .io_n_in_2(rules_42_io_n_in_2),
    .io_n_in_3(rules_42_io_n_in_3),
    .io_n_in_4(rules_42_io_n_in_4),
    .io_n_in_5(rules_42_io_n_in_5),
    .io_n_in_6(rules_42_io_n_in_6),
    .io_n_in_7(rules_42_io_n_in_7),
    .io_n_in_8(rules_42_io_n_in_8),
    .io_n_in_9(rules_42_io_n_in_9),
    .io_n_in_10(rules_42_io_n_in_10),
    .io_n_in_11(rules_42_io_n_in_11),
    .io_n_in_12(rules_42_io_n_in_12),
    .io_n_in_13(rules_42_io_n_in_13),
    .io_n_in_14(rules_42_io_n_in_14),
    .io_n_in_15(rules_42_io_n_in_15),
    .io_n_in_16(rules_42_io_n_in_16),
    .io_n_out_0(rules_42_io_n_out_0),
    .io_n_out_1(rules_42_io_n_out_1),
    .io_n_out_2(rules_42_io_n_out_2),
    .io_n_out_3(rules_42_io_n_out_3),
    .io_n_out_4(rules_42_io_n_out_4),
    .io_n_out_5(rules_42_io_n_out_5),
    .io_n_out_6(rules_42_io_n_out_6),
    .io_n_out_7(rules_42_io_n_out_7),
    .io_n_out_8(rules_42_io_n_out_8),
    .io_n_out_9(rules_42_io_n_out_9),
    .io_n_out_10(rules_42_io_n_out_10),
    .io_n_out_11(rules_42_io_n_out_11),
    .io_n_out_12(rules_42_io_n_out_12),
    .io_n_out_13(rules_42_io_n_out_13),
    .io_n_out_14(rules_42_io_n_out_14),
    .io_n_out_15(rules_42_io_n_out_15),
    .io_n_out_16(rules_42_io_n_out_16),
    .io_x_in(rules_42_io_x_in),
    .io_x_out(rules_42_io_x_out)
  );
  Exit_10 rules_43 ( // @[system.scala 24:16]
    .io_en_r(rules_43_io_en_r),
    .io_n_in_0(rules_43_io_n_in_0),
    .io_n_in_1(rules_43_io_n_in_1),
    .io_n_in_2(rules_43_io_n_in_2),
    .io_n_in_3(rules_43_io_n_in_3),
    .io_n_in_4(rules_43_io_n_in_4),
    .io_n_in_5(rules_43_io_n_in_5),
    .io_n_in_6(rules_43_io_n_in_6),
    .io_n_in_7(rules_43_io_n_in_7),
    .io_n_in_8(rules_43_io_n_in_8),
    .io_n_in_9(rules_43_io_n_in_9),
    .io_n_in_10(rules_43_io_n_in_10),
    .io_n_in_11(rules_43_io_n_in_11),
    .io_n_in_12(rules_43_io_n_in_12),
    .io_n_in_13(rules_43_io_n_in_13),
    .io_n_in_14(rules_43_io_n_in_14),
    .io_n_in_15(rules_43_io_n_in_15),
    .io_n_in_16(rules_43_io_n_in_16),
    .io_n_out_0(rules_43_io_n_out_0),
    .io_n_out_1(rules_43_io_n_out_1),
    .io_n_out_2(rules_43_io_n_out_2),
    .io_n_out_3(rules_43_io_n_out_3),
    .io_n_out_4(rules_43_io_n_out_4),
    .io_n_out_5(rules_43_io_n_out_5),
    .io_n_out_6(rules_43_io_n_out_6),
    .io_n_out_7(rules_43_io_n_out_7),
    .io_n_out_8(rules_43_io_n_out_8),
    .io_n_out_9(rules_43_io_n_out_9),
    .io_n_out_10(rules_43_io_n_out_10),
    .io_n_out_11(rules_43_io_n_out_11),
    .io_n_out_12(rules_43_io_n_out_12),
    .io_n_out_13(rules_43_io_n_out_13),
    .io_n_out_14(rules_43_io_n_out_14),
    .io_n_out_15(rules_43_io_n_out_15),
    .io_n_out_16(rules_43_io_n_out_16),
    .io_x_in(rules_43_io_x_in),
    .io_x_out(rules_43_io_x_out)
  );
  Exit_11 rules_44 ( // @[system.scala 24:16]
    .io_en_r(rules_44_io_en_r),
    .io_n_in_0(rules_44_io_n_in_0),
    .io_n_in_1(rules_44_io_n_in_1),
    .io_n_in_2(rules_44_io_n_in_2),
    .io_n_in_3(rules_44_io_n_in_3),
    .io_n_in_4(rules_44_io_n_in_4),
    .io_n_in_5(rules_44_io_n_in_5),
    .io_n_in_6(rules_44_io_n_in_6),
    .io_n_in_7(rules_44_io_n_in_7),
    .io_n_in_8(rules_44_io_n_in_8),
    .io_n_in_9(rules_44_io_n_in_9),
    .io_n_in_10(rules_44_io_n_in_10),
    .io_n_in_11(rules_44_io_n_in_11),
    .io_n_in_12(rules_44_io_n_in_12),
    .io_n_in_13(rules_44_io_n_in_13),
    .io_n_in_14(rules_44_io_n_in_14),
    .io_n_in_15(rules_44_io_n_in_15),
    .io_n_in_16(rules_44_io_n_in_16),
    .io_n_out_0(rules_44_io_n_out_0),
    .io_n_out_1(rules_44_io_n_out_1),
    .io_n_out_2(rules_44_io_n_out_2),
    .io_n_out_3(rules_44_io_n_out_3),
    .io_n_out_4(rules_44_io_n_out_4),
    .io_n_out_5(rules_44_io_n_out_5),
    .io_n_out_6(rules_44_io_n_out_6),
    .io_n_out_7(rules_44_io_n_out_7),
    .io_n_out_8(rules_44_io_n_out_8),
    .io_n_out_9(rules_44_io_n_out_9),
    .io_n_out_10(rules_44_io_n_out_10),
    .io_n_out_11(rules_44_io_n_out_11),
    .io_n_out_12(rules_44_io_n_out_12),
    .io_n_out_13(rules_44_io_n_out_13),
    .io_n_out_14(rules_44_io_n_out_14),
    .io_n_out_15(rules_44_io_n_out_15),
    .io_n_out_16(rules_44_io_n_out_16),
    .io_x_in(rules_44_io_x_in),
    .io_x_out(rules_44_io_x_out)
  );
  Exit_12 rules_45 ( // @[system.scala 24:16]
    .io_en_r(rules_45_io_en_r),
    .io_n_in_0(rules_45_io_n_in_0),
    .io_n_in_1(rules_45_io_n_in_1),
    .io_n_in_2(rules_45_io_n_in_2),
    .io_n_in_3(rules_45_io_n_in_3),
    .io_n_in_4(rules_45_io_n_in_4),
    .io_n_in_5(rules_45_io_n_in_5),
    .io_n_in_6(rules_45_io_n_in_6),
    .io_n_in_7(rules_45_io_n_in_7),
    .io_n_in_8(rules_45_io_n_in_8),
    .io_n_in_9(rules_45_io_n_in_9),
    .io_n_in_10(rules_45_io_n_in_10),
    .io_n_in_11(rules_45_io_n_in_11),
    .io_n_in_12(rules_45_io_n_in_12),
    .io_n_in_13(rules_45_io_n_in_13),
    .io_n_in_14(rules_45_io_n_in_14),
    .io_n_in_15(rules_45_io_n_in_15),
    .io_n_in_16(rules_45_io_n_in_16),
    .io_n_out_0(rules_45_io_n_out_0),
    .io_n_out_1(rules_45_io_n_out_1),
    .io_n_out_2(rules_45_io_n_out_2),
    .io_n_out_3(rules_45_io_n_out_3),
    .io_n_out_4(rules_45_io_n_out_4),
    .io_n_out_5(rules_45_io_n_out_5),
    .io_n_out_6(rules_45_io_n_out_6),
    .io_n_out_7(rules_45_io_n_out_7),
    .io_n_out_8(rules_45_io_n_out_8),
    .io_n_out_9(rules_45_io_n_out_9),
    .io_n_out_10(rules_45_io_n_out_10),
    .io_n_out_11(rules_45_io_n_out_11),
    .io_n_out_12(rules_45_io_n_out_12),
    .io_n_out_13(rules_45_io_n_out_13),
    .io_n_out_14(rules_45_io_n_out_14),
    .io_n_out_15(rules_45_io_n_out_15),
    .io_n_out_16(rules_45_io_n_out_16),
    .io_x_in(rules_45_io_x_in),
    .io_x_out(rules_45_io_x_out)
  );
  Exit_13 rules_46 ( // @[system.scala 24:16]
    .io_en_r(rules_46_io_en_r),
    .io_n_in_0(rules_46_io_n_in_0),
    .io_n_in_1(rules_46_io_n_in_1),
    .io_n_in_2(rules_46_io_n_in_2),
    .io_n_in_3(rules_46_io_n_in_3),
    .io_n_in_4(rules_46_io_n_in_4),
    .io_n_in_5(rules_46_io_n_in_5),
    .io_n_in_6(rules_46_io_n_in_6),
    .io_n_in_7(rules_46_io_n_in_7),
    .io_n_in_8(rules_46_io_n_in_8),
    .io_n_in_9(rules_46_io_n_in_9),
    .io_n_in_10(rules_46_io_n_in_10),
    .io_n_in_11(rules_46_io_n_in_11),
    .io_n_in_12(rules_46_io_n_in_12),
    .io_n_in_13(rules_46_io_n_in_13),
    .io_n_in_14(rules_46_io_n_in_14),
    .io_n_in_15(rules_46_io_n_in_15),
    .io_n_in_16(rules_46_io_n_in_16),
    .io_n_out_0(rules_46_io_n_out_0),
    .io_n_out_1(rules_46_io_n_out_1),
    .io_n_out_2(rules_46_io_n_out_2),
    .io_n_out_3(rules_46_io_n_out_3),
    .io_n_out_4(rules_46_io_n_out_4),
    .io_n_out_5(rules_46_io_n_out_5),
    .io_n_out_6(rules_46_io_n_out_6),
    .io_n_out_7(rules_46_io_n_out_7),
    .io_n_out_8(rules_46_io_n_out_8),
    .io_n_out_9(rules_46_io_n_out_9),
    .io_n_out_10(rules_46_io_n_out_10),
    .io_n_out_11(rules_46_io_n_out_11),
    .io_n_out_12(rules_46_io_n_out_12),
    .io_n_out_13(rules_46_io_n_out_13),
    .io_n_out_14(rules_46_io_n_out_14),
    .io_n_out_15(rules_46_io_n_out_15),
    .io_n_out_16(rules_46_io_n_out_16),
    .io_x_in(rules_46_io_x_in),
    .io_x_out(rules_46_io_x_out)
  );
  Exit_14 rules_47 ( // @[system.scala 24:16]
    .io_en_r(rules_47_io_en_r),
    .io_n_in_0(rules_47_io_n_in_0),
    .io_n_in_1(rules_47_io_n_in_1),
    .io_n_in_2(rules_47_io_n_in_2),
    .io_n_in_3(rules_47_io_n_in_3),
    .io_n_in_4(rules_47_io_n_in_4),
    .io_n_in_5(rules_47_io_n_in_5),
    .io_n_in_6(rules_47_io_n_in_6),
    .io_n_in_7(rules_47_io_n_in_7),
    .io_n_in_8(rules_47_io_n_in_8),
    .io_n_in_9(rules_47_io_n_in_9),
    .io_n_in_10(rules_47_io_n_in_10),
    .io_n_in_11(rules_47_io_n_in_11),
    .io_n_in_12(rules_47_io_n_in_12),
    .io_n_in_13(rules_47_io_n_in_13),
    .io_n_in_14(rules_47_io_n_in_14),
    .io_n_in_15(rules_47_io_n_in_15),
    .io_n_in_16(rules_47_io_n_in_16),
    .io_n_out_0(rules_47_io_n_out_0),
    .io_n_out_1(rules_47_io_n_out_1),
    .io_n_out_2(rules_47_io_n_out_2),
    .io_n_out_3(rules_47_io_n_out_3),
    .io_n_out_4(rules_47_io_n_out_4),
    .io_n_out_5(rules_47_io_n_out_5),
    .io_n_out_6(rules_47_io_n_out_6),
    .io_n_out_7(rules_47_io_n_out_7),
    .io_n_out_8(rules_47_io_n_out_8),
    .io_n_out_9(rules_47_io_n_out_9),
    .io_n_out_10(rules_47_io_n_out_10),
    .io_n_out_11(rules_47_io_n_out_11),
    .io_n_out_12(rules_47_io_n_out_12),
    .io_n_out_13(rules_47_io_n_out_13),
    .io_n_out_14(rules_47_io_n_out_14),
    .io_n_out_15(rules_47_io_n_out_15),
    .io_n_out_16(rules_47_io_n_out_16),
    .io_x_in(rules_47_io_x_in),
    .io_x_out(rules_47_io_x_out)
  );
  Exit_15 rules_48 ( // @[system.scala 24:16]
    .io_en_r(rules_48_io_en_r),
    .io_n_in_0(rules_48_io_n_in_0),
    .io_n_in_1(rules_48_io_n_in_1),
    .io_n_in_2(rules_48_io_n_in_2),
    .io_n_in_3(rules_48_io_n_in_3),
    .io_n_in_4(rules_48_io_n_in_4),
    .io_n_in_5(rules_48_io_n_in_5),
    .io_n_in_6(rules_48_io_n_in_6),
    .io_n_in_7(rules_48_io_n_in_7),
    .io_n_in_8(rules_48_io_n_in_8),
    .io_n_in_9(rules_48_io_n_in_9),
    .io_n_in_10(rules_48_io_n_in_10),
    .io_n_in_11(rules_48_io_n_in_11),
    .io_n_in_12(rules_48_io_n_in_12),
    .io_n_in_13(rules_48_io_n_in_13),
    .io_n_in_14(rules_48_io_n_in_14),
    .io_n_in_15(rules_48_io_n_in_15),
    .io_n_in_16(rules_48_io_n_in_16),
    .io_n_out_0(rules_48_io_n_out_0),
    .io_n_out_1(rules_48_io_n_out_1),
    .io_n_out_2(rules_48_io_n_out_2),
    .io_n_out_3(rules_48_io_n_out_3),
    .io_n_out_4(rules_48_io_n_out_4),
    .io_n_out_5(rules_48_io_n_out_5),
    .io_n_out_6(rules_48_io_n_out_6),
    .io_n_out_7(rules_48_io_n_out_7),
    .io_n_out_8(rules_48_io_n_out_8),
    .io_n_out_9(rules_48_io_n_out_9),
    .io_n_out_10(rules_48_io_n_out_10),
    .io_n_out_11(rules_48_io_n_out_11),
    .io_n_out_12(rules_48_io_n_out_12),
    .io_n_out_13(rules_48_io_n_out_13),
    .io_n_out_14(rules_48_io_n_out_14),
    .io_n_out_15(rules_48_io_n_out_15),
    .io_n_out_16(rules_48_io_n_out_16),
    .io_x_in(rules_48_io_x_in),
    .io_x_out(rules_48_io_x_out)
  );
  Idle rules_49 ( // @[system.scala 27:16]
    .io_en_r(rules_49_io_en_r),
    .io_n_in_0(rules_49_io_n_in_0),
    .io_n_in_1(rules_49_io_n_in_1),
    .io_n_in_2(rules_49_io_n_in_2),
    .io_n_in_3(rules_49_io_n_in_3),
    .io_n_in_4(rules_49_io_n_in_4),
    .io_n_in_5(rules_49_io_n_in_5),
    .io_n_in_6(rules_49_io_n_in_6),
    .io_n_in_7(rules_49_io_n_in_7),
    .io_n_in_8(rules_49_io_n_in_8),
    .io_n_in_9(rules_49_io_n_in_9),
    .io_n_in_10(rules_49_io_n_in_10),
    .io_n_in_11(rules_49_io_n_in_11),
    .io_n_in_12(rules_49_io_n_in_12),
    .io_n_in_13(rules_49_io_n_in_13),
    .io_n_in_14(rules_49_io_n_in_14),
    .io_n_in_15(rules_49_io_n_in_15),
    .io_n_in_16(rules_49_io_n_in_16),
    .io_n_out_0(rules_49_io_n_out_0),
    .io_n_out_1(rules_49_io_n_out_1),
    .io_n_out_2(rules_49_io_n_out_2),
    .io_n_out_3(rules_49_io_n_out_3),
    .io_n_out_4(rules_49_io_n_out_4),
    .io_n_out_5(rules_49_io_n_out_5),
    .io_n_out_6(rules_49_io_n_out_6),
    .io_n_out_7(rules_49_io_n_out_7),
    .io_n_out_8(rules_49_io_n_out_8),
    .io_n_out_9(rules_49_io_n_out_9),
    .io_n_out_10(rules_49_io_n_out_10),
    .io_n_out_11(rules_49_io_n_out_11),
    .io_n_out_12(rules_49_io_n_out_12),
    .io_n_out_13(rules_49_io_n_out_13),
    .io_n_out_14(rules_49_io_n_out_14),
    .io_n_out_15(rules_49_io_n_out_15),
    .io_n_out_16(rules_49_io_n_out_16),
    .io_x_in(rules_49_io_x_in),
    .io_x_out(rules_49_io_x_out)
  );
  Idle_1 rules_50 ( // @[system.scala 27:16]
    .io_en_r(rules_50_io_en_r),
    .io_n_in_0(rules_50_io_n_in_0),
    .io_n_in_1(rules_50_io_n_in_1),
    .io_n_in_2(rules_50_io_n_in_2),
    .io_n_in_3(rules_50_io_n_in_3),
    .io_n_in_4(rules_50_io_n_in_4),
    .io_n_in_5(rules_50_io_n_in_5),
    .io_n_in_6(rules_50_io_n_in_6),
    .io_n_in_7(rules_50_io_n_in_7),
    .io_n_in_8(rules_50_io_n_in_8),
    .io_n_in_9(rules_50_io_n_in_9),
    .io_n_in_10(rules_50_io_n_in_10),
    .io_n_in_11(rules_50_io_n_in_11),
    .io_n_in_12(rules_50_io_n_in_12),
    .io_n_in_13(rules_50_io_n_in_13),
    .io_n_in_14(rules_50_io_n_in_14),
    .io_n_in_15(rules_50_io_n_in_15),
    .io_n_in_16(rules_50_io_n_in_16),
    .io_n_out_0(rules_50_io_n_out_0),
    .io_n_out_1(rules_50_io_n_out_1),
    .io_n_out_2(rules_50_io_n_out_2),
    .io_n_out_3(rules_50_io_n_out_3),
    .io_n_out_4(rules_50_io_n_out_4),
    .io_n_out_5(rules_50_io_n_out_5),
    .io_n_out_6(rules_50_io_n_out_6),
    .io_n_out_7(rules_50_io_n_out_7),
    .io_n_out_8(rules_50_io_n_out_8),
    .io_n_out_9(rules_50_io_n_out_9),
    .io_n_out_10(rules_50_io_n_out_10),
    .io_n_out_11(rules_50_io_n_out_11),
    .io_n_out_12(rules_50_io_n_out_12),
    .io_n_out_13(rules_50_io_n_out_13),
    .io_n_out_14(rules_50_io_n_out_14),
    .io_n_out_15(rules_50_io_n_out_15),
    .io_n_out_16(rules_50_io_n_out_16),
    .io_x_in(rules_50_io_x_in),
    .io_x_out(rules_50_io_x_out)
  );
  Idle_2 rules_51 ( // @[system.scala 27:16]
    .io_en_r(rules_51_io_en_r),
    .io_n_in_0(rules_51_io_n_in_0),
    .io_n_in_1(rules_51_io_n_in_1),
    .io_n_in_2(rules_51_io_n_in_2),
    .io_n_in_3(rules_51_io_n_in_3),
    .io_n_in_4(rules_51_io_n_in_4),
    .io_n_in_5(rules_51_io_n_in_5),
    .io_n_in_6(rules_51_io_n_in_6),
    .io_n_in_7(rules_51_io_n_in_7),
    .io_n_in_8(rules_51_io_n_in_8),
    .io_n_in_9(rules_51_io_n_in_9),
    .io_n_in_10(rules_51_io_n_in_10),
    .io_n_in_11(rules_51_io_n_in_11),
    .io_n_in_12(rules_51_io_n_in_12),
    .io_n_in_13(rules_51_io_n_in_13),
    .io_n_in_14(rules_51_io_n_in_14),
    .io_n_in_15(rules_51_io_n_in_15),
    .io_n_in_16(rules_51_io_n_in_16),
    .io_n_out_0(rules_51_io_n_out_0),
    .io_n_out_1(rules_51_io_n_out_1),
    .io_n_out_2(rules_51_io_n_out_2),
    .io_n_out_3(rules_51_io_n_out_3),
    .io_n_out_4(rules_51_io_n_out_4),
    .io_n_out_5(rules_51_io_n_out_5),
    .io_n_out_6(rules_51_io_n_out_6),
    .io_n_out_7(rules_51_io_n_out_7),
    .io_n_out_8(rules_51_io_n_out_8),
    .io_n_out_9(rules_51_io_n_out_9),
    .io_n_out_10(rules_51_io_n_out_10),
    .io_n_out_11(rules_51_io_n_out_11),
    .io_n_out_12(rules_51_io_n_out_12),
    .io_n_out_13(rules_51_io_n_out_13),
    .io_n_out_14(rules_51_io_n_out_14),
    .io_n_out_15(rules_51_io_n_out_15),
    .io_n_out_16(rules_51_io_n_out_16),
    .io_x_in(rules_51_io_x_in),
    .io_x_out(rules_51_io_x_out)
  );
  Idle_3 rules_52 ( // @[system.scala 27:16]
    .io_en_r(rules_52_io_en_r),
    .io_n_in_0(rules_52_io_n_in_0),
    .io_n_in_1(rules_52_io_n_in_1),
    .io_n_in_2(rules_52_io_n_in_2),
    .io_n_in_3(rules_52_io_n_in_3),
    .io_n_in_4(rules_52_io_n_in_4),
    .io_n_in_5(rules_52_io_n_in_5),
    .io_n_in_6(rules_52_io_n_in_6),
    .io_n_in_7(rules_52_io_n_in_7),
    .io_n_in_8(rules_52_io_n_in_8),
    .io_n_in_9(rules_52_io_n_in_9),
    .io_n_in_10(rules_52_io_n_in_10),
    .io_n_in_11(rules_52_io_n_in_11),
    .io_n_in_12(rules_52_io_n_in_12),
    .io_n_in_13(rules_52_io_n_in_13),
    .io_n_in_14(rules_52_io_n_in_14),
    .io_n_in_15(rules_52_io_n_in_15),
    .io_n_in_16(rules_52_io_n_in_16),
    .io_n_out_0(rules_52_io_n_out_0),
    .io_n_out_1(rules_52_io_n_out_1),
    .io_n_out_2(rules_52_io_n_out_2),
    .io_n_out_3(rules_52_io_n_out_3),
    .io_n_out_4(rules_52_io_n_out_4),
    .io_n_out_5(rules_52_io_n_out_5),
    .io_n_out_6(rules_52_io_n_out_6),
    .io_n_out_7(rules_52_io_n_out_7),
    .io_n_out_8(rules_52_io_n_out_8),
    .io_n_out_9(rules_52_io_n_out_9),
    .io_n_out_10(rules_52_io_n_out_10),
    .io_n_out_11(rules_52_io_n_out_11),
    .io_n_out_12(rules_52_io_n_out_12),
    .io_n_out_13(rules_52_io_n_out_13),
    .io_n_out_14(rules_52_io_n_out_14),
    .io_n_out_15(rules_52_io_n_out_15),
    .io_n_out_16(rules_52_io_n_out_16),
    .io_x_in(rules_52_io_x_in),
    .io_x_out(rules_52_io_x_out)
  );
  Idle_4 rules_53 ( // @[system.scala 27:16]
    .io_en_r(rules_53_io_en_r),
    .io_n_in_0(rules_53_io_n_in_0),
    .io_n_in_1(rules_53_io_n_in_1),
    .io_n_in_2(rules_53_io_n_in_2),
    .io_n_in_3(rules_53_io_n_in_3),
    .io_n_in_4(rules_53_io_n_in_4),
    .io_n_in_5(rules_53_io_n_in_5),
    .io_n_in_6(rules_53_io_n_in_6),
    .io_n_in_7(rules_53_io_n_in_7),
    .io_n_in_8(rules_53_io_n_in_8),
    .io_n_in_9(rules_53_io_n_in_9),
    .io_n_in_10(rules_53_io_n_in_10),
    .io_n_in_11(rules_53_io_n_in_11),
    .io_n_in_12(rules_53_io_n_in_12),
    .io_n_in_13(rules_53_io_n_in_13),
    .io_n_in_14(rules_53_io_n_in_14),
    .io_n_in_15(rules_53_io_n_in_15),
    .io_n_in_16(rules_53_io_n_in_16),
    .io_n_out_0(rules_53_io_n_out_0),
    .io_n_out_1(rules_53_io_n_out_1),
    .io_n_out_2(rules_53_io_n_out_2),
    .io_n_out_3(rules_53_io_n_out_3),
    .io_n_out_4(rules_53_io_n_out_4),
    .io_n_out_5(rules_53_io_n_out_5),
    .io_n_out_6(rules_53_io_n_out_6),
    .io_n_out_7(rules_53_io_n_out_7),
    .io_n_out_8(rules_53_io_n_out_8),
    .io_n_out_9(rules_53_io_n_out_9),
    .io_n_out_10(rules_53_io_n_out_10),
    .io_n_out_11(rules_53_io_n_out_11),
    .io_n_out_12(rules_53_io_n_out_12),
    .io_n_out_13(rules_53_io_n_out_13),
    .io_n_out_14(rules_53_io_n_out_14),
    .io_n_out_15(rules_53_io_n_out_15),
    .io_n_out_16(rules_53_io_n_out_16),
    .io_x_in(rules_53_io_x_in),
    .io_x_out(rules_53_io_x_out)
  );
  Idle_5 rules_54 ( // @[system.scala 27:16]
    .io_en_r(rules_54_io_en_r),
    .io_n_in_0(rules_54_io_n_in_0),
    .io_n_in_1(rules_54_io_n_in_1),
    .io_n_in_2(rules_54_io_n_in_2),
    .io_n_in_3(rules_54_io_n_in_3),
    .io_n_in_4(rules_54_io_n_in_4),
    .io_n_in_5(rules_54_io_n_in_5),
    .io_n_in_6(rules_54_io_n_in_6),
    .io_n_in_7(rules_54_io_n_in_7),
    .io_n_in_8(rules_54_io_n_in_8),
    .io_n_in_9(rules_54_io_n_in_9),
    .io_n_in_10(rules_54_io_n_in_10),
    .io_n_in_11(rules_54_io_n_in_11),
    .io_n_in_12(rules_54_io_n_in_12),
    .io_n_in_13(rules_54_io_n_in_13),
    .io_n_in_14(rules_54_io_n_in_14),
    .io_n_in_15(rules_54_io_n_in_15),
    .io_n_in_16(rules_54_io_n_in_16),
    .io_n_out_0(rules_54_io_n_out_0),
    .io_n_out_1(rules_54_io_n_out_1),
    .io_n_out_2(rules_54_io_n_out_2),
    .io_n_out_3(rules_54_io_n_out_3),
    .io_n_out_4(rules_54_io_n_out_4),
    .io_n_out_5(rules_54_io_n_out_5),
    .io_n_out_6(rules_54_io_n_out_6),
    .io_n_out_7(rules_54_io_n_out_7),
    .io_n_out_8(rules_54_io_n_out_8),
    .io_n_out_9(rules_54_io_n_out_9),
    .io_n_out_10(rules_54_io_n_out_10),
    .io_n_out_11(rules_54_io_n_out_11),
    .io_n_out_12(rules_54_io_n_out_12),
    .io_n_out_13(rules_54_io_n_out_13),
    .io_n_out_14(rules_54_io_n_out_14),
    .io_n_out_15(rules_54_io_n_out_15),
    .io_n_out_16(rules_54_io_n_out_16),
    .io_x_in(rules_54_io_x_in),
    .io_x_out(rules_54_io_x_out)
  );
  Idle_6 rules_55 ( // @[system.scala 27:16]
    .io_en_r(rules_55_io_en_r),
    .io_n_in_0(rules_55_io_n_in_0),
    .io_n_in_1(rules_55_io_n_in_1),
    .io_n_in_2(rules_55_io_n_in_2),
    .io_n_in_3(rules_55_io_n_in_3),
    .io_n_in_4(rules_55_io_n_in_4),
    .io_n_in_5(rules_55_io_n_in_5),
    .io_n_in_6(rules_55_io_n_in_6),
    .io_n_in_7(rules_55_io_n_in_7),
    .io_n_in_8(rules_55_io_n_in_8),
    .io_n_in_9(rules_55_io_n_in_9),
    .io_n_in_10(rules_55_io_n_in_10),
    .io_n_in_11(rules_55_io_n_in_11),
    .io_n_in_12(rules_55_io_n_in_12),
    .io_n_in_13(rules_55_io_n_in_13),
    .io_n_in_14(rules_55_io_n_in_14),
    .io_n_in_15(rules_55_io_n_in_15),
    .io_n_in_16(rules_55_io_n_in_16),
    .io_n_out_0(rules_55_io_n_out_0),
    .io_n_out_1(rules_55_io_n_out_1),
    .io_n_out_2(rules_55_io_n_out_2),
    .io_n_out_3(rules_55_io_n_out_3),
    .io_n_out_4(rules_55_io_n_out_4),
    .io_n_out_5(rules_55_io_n_out_5),
    .io_n_out_6(rules_55_io_n_out_6),
    .io_n_out_7(rules_55_io_n_out_7),
    .io_n_out_8(rules_55_io_n_out_8),
    .io_n_out_9(rules_55_io_n_out_9),
    .io_n_out_10(rules_55_io_n_out_10),
    .io_n_out_11(rules_55_io_n_out_11),
    .io_n_out_12(rules_55_io_n_out_12),
    .io_n_out_13(rules_55_io_n_out_13),
    .io_n_out_14(rules_55_io_n_out_14),
    .io_n_out_15(rules_55_io_n_out_15),
    .io_n_out_16(rules_55_io_n_out_16),
    .io_x_in(rules_55_io_x_in),
    .io_x_out(rules_55_io_x_out)
  );
  Idle_7 rules_56 ( // @[system.scala 27:16]
    .io_en_r(rules_56_io_en_r),
    .io_n_in_0(rules_56_io_n_in_0),
    .io_n_in_1(rules_56_io_n_in_1),
    .io_n_in_2(rules_56_io_n_in_2),
    .io_n_in_3(rules_56_io_n_in_3),
    .io_n_in_4(rules_56_io_n_in_4),
    .io_n_in_5(rules_56_io_n_in_5),
    .io_n_in_6(rules_56_io_n_in_6),
    .io_n_in_7(rules_56_io_n_in_7),
    .io_n_in_8(rules_56_io_n_in_8),
    .io_n_in_9(rules_56_io_n_in_9),
    .io_n_in_10(rules_56_io_n_in_10),
    .io_n_in_11(rules_56_io_n_in_11),
    .io_n_in_12(rules_56_io_n_in_12),
    .io_n_in_13(rules_56_io_n_in_13),
    .io_n_in_14(rules_56_io_n_in_14),
    .io_n_in_15(rules_56_io_n_in_15),
    .io_n_in_16(rules_56_io_n_in_16),
    .io_n_out_0(rules_56_io_n_out_0),
    .io_n_out_1(rules_56_io_n_out_1),
    .io_n_out_2(rules_56_io_n_out_2),
    .io_n_out_3(rules_56_io_n_out_3),
    .io_n_out_4(rules_56_io_n_out_4),
    .io_n_out_5(rules_56_io_n_out_5),
    .io_n_out_6(rules_56_io_n_out_6),
    .io_n_out_7(rules_56_io_n_out_7),
    .io_n_out_8(rules_56_io_n_out_8),
    .io_n_out_9(rules_56_io_n_out_9),
    .io_n_out_10(rules_56_io_n_out_10),
    .io_n_out_11(rules_56_io_n_out_11),
    .io_n_out_12(rules_56_io_n_out_12),
    .io_n_out_13(rules_56_io_n_out_13),
    .io_n_out_14(rules_56_io_n_out_14),
    .io_n_out_15(rules_56_io_n_out_15),
    .io_n_out_16(rules_56_io_n_out_16),
    .io_x_in(rules_56_io_x_in),
    .io_x_out(rules_56_io_x_out)
  );
  Idle_8 rules_57 ( // @[system.scala 27:16]
    .io_en_r(rules_57_io_en_r),
    .io_n_in_0(rules_57_io_n_in_0),
    .io_n_in_1(rules_57_io_n_in_1),
    .io_n_in_2(rules_57_io_n_in_2),
    .io_n_in_3(rules_57_io_n_in_3),
    .io_n_in_4(rules_57_io_n_in_4),
    .io_n_in_5(rules_57_io_n_in_5),
    .io_n_in_6(rules_57_io_n_in_6),
    .io_n_in_7(rules_57_io_n_in_7),
    .io_n_in_8(rules_57_io_n_in_8),
    .io_n_in_9(rules_57_io_n_in_9),
    .io_n_in_10(rules_57_io_n_in_10),
    .io_n_in_11(rules_57_io_n_in_11),
    .io_n_in_12(rules_57_io_n_in_12),
    .io_n_in_13(rules_57_io_n_in_13),
    .io_n_in_14(rules_57_io_n_in_14),
    .io_n_in_15(rules_57_io_n_in_15),
    .io_n_in_16(rules_57_io_n_in_16),
    .io_n_out_0(rules_57_io_n_out_0),
    .io_n_out_1(rules_57_io_n_out_1),
    .io_n_out_2(rules_57_io_n_out_2),
    .io_n_out_3(rules_57_io_n_out_3),
    .io_n_out_4(rules_57_io_n_out_4),
    .io_n_out_5(rules_57_io_n_out_5),
    .io_n_out_6(rules_57_io_n_out_6),
    .io_n_out_7(rules_57_io_n_out_7),
    .io_n_out_8(rules_57_io_n_out_8),
    .io_n_out_9(rules_57_io_n_out_9),
    .io_n_out_10(rules_57_io_n_out_10),
    .io_n_out_11(rules_57_io_n_out_11),
    .io_n_out_12(rules_57_io_n_out_12),
    .io_n_out_13(rules_57_io_n_out_13),
    .io_n_out_14(rules_57_io_n_out_14),
    .io_n_out_15(rules_57_io_n_out_15),
    .io_n_out_16(rules_57_io_n_out_16),
    .io_x_in(rules_57_io_x_in),
    .io_x_out(rules_57_io_x_out)
  );
  Idle_9 rules_58 ( // @[system.scala 27:16]
    .io_en_r(rules_58_io_en_r),
    .io_n_in_0(rules_58_io_n_in_0),
    .io_n_in_1(rules_58_io_n_in_1),
    .io_n_in_2(rules_58_io_n_in_2),
    .io_n_in_3(rules_58_io_n_in_3),
    .io_n_in_4(rules_58_io_n_in_4),
    .io_n_in_5(rules_58_io_n_in_5),
    .io_n_in_6(rules_58_io_n_in_6),
    .io_n_in_7(rules_58_io_n_in_7),
    .io_n_in_8(rules_58_io_n_in_8),
    .io_n_in_9(rules_58_io_n_in_9),
    .io_n_in_10(rules_58_io_n_in_10),
    .io_n_in_11(rules_58_io_n_in_11),
    .io_n_in_12(rules_58_io_n_in_12),
    .io_n_in_13(rules_58_io_n_in_13),
    .io_n_in_14(rules_58_io_n_in_14),
    .io_n_in_15(rules_58_io_n_in_15),
    .io_n_in_16(rules_58_io_n_in_16),
    .io_n_out_0(rules_58_io_n_out_0),
    .io_n_out_1(rules_58_io_n_out_1),
    .io_n_out_2(rules_58_io_n_out_2),
    .io_n_out_3(rules_58_io_n_out_3),
    .io_n_out_4(rules_58_io_n_out_4),
    .io_n_out_5(rules_58_io_n_out_5),
    .io_n_out_6(rules_58_io_n_out_6),
    .io_n_out_7(rules_58_io_n_out_7),
    .io_n_out_8(rules_58_io_n_out_8),
    .io_n_out_9(rules_58_io_n_out_9),
    .io_n_out_10(rules_58_io_n_out_10),
    .io_n_out_11(rules_58_io_n_out_11),
    .io_n_out_12(rules_58_io_n_out_12),
    .io_n_out_13(rules_58_io_n_out_13),
    .io_n_out_14(rules_58_io_n_out_14),
    .io_n_out_15(rules_58_io_n_out_15),
    .io_n_out_16(rules_58_io_n_out_16),
    .io_x_in(rules_58_io_x_in),
    .io_x_out(rules_58_io_x_out)
  );
  Idle_10 rules_59 ( // @[system.scala 27:16]
    .io_en_r(rules_59_io_en_r),
    .io_n_in_0(rules_59_io_n_in_0),
    .io_n_in_1(rules_59_io_n_in_1),
    .io_n_in_2(rules_59_io_n_in_2),
    .io_n_in_3(rules_59_io_n_in_3),
    .io_n_in_4(rules_59_io_n_in_4),
    .io_n_in_5(rules_59_io_n_in_5),
    .io_n_in_6(rules_59_io_n_in_6),
    .io_n_in_7(rules_59_io_n_in_7),
    .io_n_in_8(rules_59_io_n_in_8),
    .io_n_in_9(rules_59_io_n_in_9),
    .io_n_in_10(rules_59_io_n_in_10),
    .io_n_in_11(rules_59_io_n_in_11),
    .io_n_in_12(rules_59_io_n_in_12),
    .io_n_in_13(rules_59_io_n_in_13),
    .io_n_in_14(rules_59_io_n_in_14),
    .io_n_in_15(rules_59_io_n_in_15),
    .io_n_in_16(rules_59_io_n_in_16),
    .io_n_out_0(rules_59_io_n_out_0),
    .io_n_out_1(rules_59_io_n_out_1),
    .io_n_out_2(rules_59_io_n_out_2),
    .io_n_out_3(rules_59_io_n_out_3),
    .io_n_out_4(rules_59_io_n_out_4),
    .io_n_out_5(rules_59_io_n_out_5),
    .io_n_out_6(rules_59_io_n_out_6),
    .io_n_out_7(rules_59_io_n_out_7),
    .io_n_out_8(rules_59_io_n_out_8),
    .io_n_out_9(rules_59_io_n_out_9),
    .io_n_out_10(rules_59_io_n_out_10),
    .io_n_out_11(rules_59_io_n_out_11),
    .io_n_out_12(rules_59_io_n_out_12),
    .io_n_out_13(rules_59_io_n_out_13),
    .io_n_out_14(rules_59_io_n_out_14),
    .io_n_out_15(rules_59_io_n_out_15),
    .io_n_out_16(rules_59_io_n_out_16),
    .io_x_in(rules_59_io_x_in),
    .io_x_out(rules_59_io_x_out)
  );
  Idle_11 rules_60 ( // @[system.scala 27:16]
    .io_en_r(rules_60_io_en_r),
    .io_n_in_0(rules_60_io_n_in_0),
    .io_n_in_1(rules_60_io_n_in_1),
    .io_n_in_2(rules_60_io_n_in_2),
    .io_n_in_3(rules_60_io_n_in_3),
    .io_n_in_4(rules_60_io_n_in_4),
    .io_n_in_5(rules_60_io_n_in_5),
    .io_n_in_6(rules_60_io_n_in_6),
    .io_n_in_7(rules_60_io_n_in_7),
    .io_n_in_8(rules_60_io_n_in_8),
    .io_n_in_9(rules_60_io_n_in_9),
    .io_n_in_10(rules_60_io_n_in_10),
    .io_n_in_11(rules_60_io_n_in_11),
    .io_n_in_12(rules_60_io_n_in_12),
    .io_n_in_13(rules_60_io_n_in_13),
    .io_n_in_14(rules_60_io_n_in_14),
    .io_n_in_15(rules_60_io_n_in_15),
    .io_n_in_16(rules_60_io_n_in_16),
    .io_n_out_0(rules_60_io_n_out_0),
    .io_n_out_1(rules_60_io_n_out_1),
    .io_n_out_2(rules_60_io_n_out_2),
    .io_n_out_3(rules_60_io_n_out_3),
    .io_n_out_4(rules_60_io_n_out_4),
    .io_n_out_5(rules_60_io_n_out_5),
    .io_n_out_6(rules_60_io_n_out_6),
    .io_n_out_7(rules_60_io_n_out_7),
    .io_n_out_8(rules_60_io_n_out_8),
    .io_n_out_9(rules_60_io_n_out_9),
    .io_n_out_10(rules_60_io_n_out_10),
    .io_n_out_11(rules_60_io_n_out_11),
    .io_n_out_12(rules_60_io_n_out_12),
    .io_n_out_13(rules_60_io_n_out_13),
    .io_n_out_14(rules_60_io_n_out_14),
    .io_n_out_15(rules_60_io_n_out_15),
    .io_n_out_16(rules_60_io_n_out_16),
    .io_x_in(rules_60_io_x_in),
    .io_x_out(rules_60_io_x_out)
  );
  Idle_12 rules_61 ( // @[system.scala 27:16]
    .io_en_r(rules_61_io_en_r),
    .io_n_in_0(rules_61_io_n_in_0),
    .io_n_in_1(rules_61_io_n_in_1),
    .io_n_in_2(rules_61_io_n_in_2),
    .io_n_in_3(rules_61_io_n_in_3),
    .io_n_in_4(rules_61_io_n_in_4),
    .io_n_in_5(rules_61_io_n_in_5),
    .io_n_in_6(rules_61_io_n_in_6),
    .io_n_in_7(rules_61_io_n_in_7),
    .io_n_in_8(rules_61_io_n_in_8),
    .io_n_in_9(rules_61_io_n_in_9),
    .io_n_in_10(rules_61_io_n_in_10),
    .io_n_in_11(rules_61_io_n_in_11),
    .io_n_in_12(rules_61_io_n_in_12),
    .io_n_in_13(rules_61_io_n_in_13),
    .io_n_in_14(rules_61_io_n_in_14),
    .io_n_in_15(rules_61_io_n_in_15),
    .io_n_in_16(rules_61_io_n_in_16),
    .io_n_out_0(rules_61_io_n_out_0),
    .io_n_out_1(rules_61_io_n_out_1),
    .io_n_out_2(rules_61_io_n_out_2),
    .io_n_out_3(rules_61_io_n_out_3),
    .io_n_out_4(rules_61_io_n_out_4),
    .io_n_out_5(rules_61_io_n_out_5),
    .io_n_out_6(rules_61_io_n_out_6),
    .io_n_out_7(rules_61_io_n_out_7),
    .io_n_out_8(rules_61_io_n_out_8),
    .io_n_out_9(rules_61_io_n_out_9),
    .io_n_out_10(rules_61_io_n_out_10),
    .io_n_out_11(rules_61_io_n_out_11),
    .io_n_out_12(rules_61_io_n_out_12),
    .io_n_out_13(rules_61_io_n_out_13),
    .io_n_out_14(rules_61_io_n_out_14),
    .io_n_out_15(rules_61_io_n_out_15),
    .io_n_out_16(rules_61_io_n_out_16),
    .io_x_in(rules_61_io_x_in),
    .io_x_out(rules_61_io_x_out)
  );
  Idle_13 rules_62 ( // @[system.scala 27:16]
    .io_en_r(rules_62_io_en_r),
    .io_n_in_0(rules_62_io_n_in_0),
    .io_n_in_1(rules_62_io_n_in_1),
    .io_n_in_2(rules_62_io_n_in_2),
    .io_n_in_3(rules_62_io_n_in_3),
    .io_n_in_4(rules_62_io_n_in_4),
    .io_n_in_5(rules_62_io_n_in_5),
    .io_n_in_6(rules_62_io_n_in_6),
    .io_n_in_7(rules_62_io_n_in_7),
    .io_n_in_8(rules_62_io_n_in_8),
    .io_n_in_9(rules_62_io_n_in_9),
    .io_n_in_10(rules_62_io_n_in_10),
    .io_n_in_11(rules_62_io_n_in_11),
    .io_n_in_12(rules_62_io_n_in_12),
    .io_n_in_13(rules_62_io_n_in_13),
    .io_n_in_14(rules_62_io_n_in_14),
    .io_n_in_15(rules_62_io_n_in_15),
    .io_n_in_16(rules_62_io_n_in_16),
    .io_n_out_0(rules_62_io_n_out_0),
    .io_n_out_1(rules_62_io_n_out_1),
    .io_n_out_2(rules_62_io_n_out_2),
    .io_n_out_3(rules_62_io_n_out_3),
    .io_n_out_4(rules_62_io_n_out_4),
    .io_n_out_5(rules_62_io_n_out_5),
    .io_n_out_6(rules_62_io_n_out_6),
    .io_n_out_7(rules_62_io_n_out_7),
    .io_n_out_8(rules_62_io_n_out_8),
    .io_n_out_9(rules_62_io_n_out_9),
    .io_n_out_10(rules_62_io_n_out_10),
    .io_n_out_11(rules_62_io_n_out_11),
    .io_n_out_12(rules_62_io_n_out_12),
    .io_n_out_13(rules_62_io_n_out_13),
    .io_n_out_14(rules_62_io_n_out_14),
    .io_n_out_15(rules_62_io_n_out_15),
    .io_n_out_16(rules_62_io_n_out_16),
    .io_x_in(rules_62_io_x_in),
    .io_x_out(rules_62_io_x_out)
  );
  Idle_14 rules_63 ( // @[system.scala 27:16]
    .io_en_r(rules_63_io_en_r),
    .io_n_in_0(rules_63_io_n_in_0),
    .io_n_in_1(rules_63_io_n_in_1),
    .io_n_in_2(rules_63_io_n_in_2),
    .io_n_in_3(rules_63_io_n_in_3),
    .io_n_in_4(rules_63_io_n_in_4),
    .io_n_in_5(rules_63_io_n_in_5),
    .io_n_in_6(rules_63_io_n_in_6),
    .io_n_in_7(rules_63_io_n_in_7),
    .io_n_in_8(rules_63_io_n_in_8),
    .io_n_in_9(rules_63_io_n_in_9),
    .io_n_in_10(rules_63_io_n_in_10),
    .io_n_in_11(rules_63_io_n_in_11),
    .io_n_in_12(rules_63_io_n_in_12),
    .io_n_in_13(rules_63_io_n_in_13),
    .io_n_in_14(rules_63_io_n_in_14),
    .io_n_in_15(rules_63_io_n_in_15),
    .io_n_in_16(rules_63_io_n_in_16),
    .io_n_out_0(rules_63_io_n_out_0),
    .io_n_out_1(rules_63_io_n_out_1),
    .io_n_out_2(rules_63_io_n_out_2),
    .io_n_out_3(rules_63_io_n_out_3),
    .io_n_out_4(rules_63_io_n_out_4),
    .io_n_out_5(rules_63_io_n_out_5),
    .io_n_out_6(rules_63_io_n_out_6),
    .io_n_out_7(rules_63_io_n_out_7),
    .io_n_out_8(rules_63_io_n_out_8),
    .io_n_out_9(rules_63_io_n_out_9),
    .io_n_out_10(rules_63_io_n_out_10),
    .io_n_out_11(rules_63_io_n_out_11),
    .io_n_out_12(rules_63_io_n_out_12),
    .io_n_out_13(rules_63_io_n_out_13),
    .io_n_out_14(rules_63_io_n_out_14),
    .io_n_out_15(rules_63_io_n_out_15),
    .io_n_out_16(rules_63_io_n_out_16),
    .io_x_in(rules_63_io_x_in),
    .io_x_out(rules_63_io_x_out)
  );
  Idle_15 rules_64 ( // @[system.scala 27:16]
    .io_en_r(rules_64_io_en_r),
    .io_n_in_0(rules_64_io_n_in_0),
    .io_n_in_1(rules_64_io_n_in_1),
    .io_n_in_2(rules_64_io_n_in_2),
    .io_n_in_3(rules_64_io_n_in_3),
    .io_n_in_4(rules_64_io_n_in_4),
    .io_n_in_5(rules_64_io_n_in_5),
    .io_n_in_6(rules_64_io_n_in_6),
    .io_n_in_7(rules_64_io_n_in_7),
    .io_n_in_8(rules_64_io_n_in_8),
    .io_n_in_9(rules_64_io_n_in_9),
    .io_n_in_10(rules_64_io_n_in_10),
    .io_n_in_11(rules_64_io_n_in_11),
    .io_n_in_12(rules_64_io_n_in_12),
    .io_n_in_13(rules_64_io_n_in_13),
    .io_n_in_14(rules_64_io_n_in_14),
    .io_n_in_15(rules_64_io_n_in_15),
    .io_n_in_16(rules_64_io_n_in_16),
    .io_n_out_0(rules_64_io_n_out_0),
    .io_n_out_1(rules_64_io_n_out_1),
    .io_n_out_2(rules_64_io_n_out_2),
    .io_n_out_3(rules_64_io_n_out_3),
    .io_n_out_4(rules_64_io_n_out_4),
    .io_n_out_5(rules_64_io_n_out_5),
    .io_n_out_6(rules_64_io_n_out_6),
    .io_n_out_7(rules_64_io_n_out_7),
    .io_n_out_8(rules_64_io_n_out_8),
    .io_n_out_9(rules_64_io_n_out_9),
    .io_n_out_10(rules_64_io_n_out_10),
    .io_n_out_11(rules_64_io_n_out_11),
    .io_n_out_12(rules_64_io_n_out_12),
    .io_n_out_13(rules_64_io_n_out_13),
    .io_n_out_14(rules_64_io_n_out_14),
    .io_n_out_15(rules_64_io_n_out_15),
    .io_n_out_16(rules_64_io_n_out_16),
    .io_x_in(rules_64_io_x_in),
    .io_x_out(rules_64_io_x_out)
  );
  assign io_n_out_0 = n_reg_0; // @[system.scala 13:9]
  assign io_n_out_1 = n_reg_1; // @[system.scala 13:9]
  assign io_n_out_2 = n_reg_2; // @[system.scala 13:9]
  assign io_n_out_3 = n_reg_3; // @[system.scala 13:9]
  assign io_n_out_4 = n_reg_4; // @[system.scala 13:9]
  assign io_n_out_5 = n_reg_5; // @[system.scala 13:9]
  assign io_n_out_6 = n_reg_6; // @[system.scala 13:9]
  assign io_n_out_7 = n_reg_7; // @[system.scala 13:9]
  assign io_n_out_8 = n_reg_8; // @[system.scala 13:9]
  assign io_n_out_9 = n_reg_9; // @[system.scala 13:9]
  assign io_n_out_10 = n_reg_10; // @[system.scala 13:9]
  assign io_n_out_11 = n_reg_11; // @[system.scala 13:9]
  assign io_n_out_12 = n_reg_12; // @[system.scala 13:9]
  assign io_n_out_13 = n_reg_13; // @[system.scala 13:9]
  assign io_n_out_14 = n_reg_14; // @[system.scala 13:9]
  assign io_n_out_15 = n_reg_15; // @[system.scala 13:9]
  assign io_n_out_16 = n_reg_16; // @[system.scala 13:9]
  assign io_x_out = x_reg; // @[system.scala 15:9]
  assign rules_0_io_en_r = io_en_a == 7'h0; // @[system.scala 32:27]
  assign rules_0_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_0_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_0_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_0_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_0_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_0_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_0_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_0_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_0_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_0_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_0_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_0_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_0_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_0_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_0_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_0_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_0_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_0_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_1_io_en_r = io_en_a == 7'h1; // @[system.scala 32:27]
  assign rules_1_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_1_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_1_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_1_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_1_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_1_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_1_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_1_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_1_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_1_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_1_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_1_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_1_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_1_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_1_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_1_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_1_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_1_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_2_io_en_r = io_en_a == 7'h2; // @[system.scala 32:27]
  assign rules_2_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_2_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_2_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_2_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_2_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_2_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_2_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_2_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_2_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_2_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_2_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_2_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_2_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_2_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_2_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_2_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_2_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_2_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_3_io_en_r = io_en_a == 7'h3; // @[system.scala 32:27]
  assign rules_3_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_3_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_3_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_3_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_3_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_3_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_3_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_3_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_3_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_3_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_3_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_3_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_3_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_3_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_3_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_3_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_3_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_3_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_4_io_en_r = io_en_a == 7'h4; // @[system.scala 32:27]
  assign rules_4_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_4_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_4_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_4_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_4_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_4_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_4_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_4_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_4_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_4_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_4_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_4_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_4_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_4_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_4_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_4_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_4_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_4_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_5_io_en_r = io_en_a == 7'h5; // @[system.scala 32:27]
  assign rules_5_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_5_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_5_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_5_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_5_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_5_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_5_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_5_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_5_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_5_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_5_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_5_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_5_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_5_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_5_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_5_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_5_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_5_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_6_io_en_r = io_en_a == 7'h6; // @[system.scala 32:27]
  assign rules_6_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_6_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_6_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_6_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_6_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_6_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_6_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_6_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_6_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_6_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_6_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_6_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_6_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_6_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_6_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_6_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_6_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_6_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_7_io_en_r = io_en_a == 7'h7; // @[system.scala 32:27]
  assign rules_7_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_7_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_7_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_7_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_7_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_7_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_7_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_7_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_7_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_7_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_7_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_7_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_7_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_7_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_7_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_7_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_7_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_7_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_8_io_en_r = io_en_a == 7'h8; // @[system.scala 32:27]
  assign rules_8_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_8_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_8_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_8_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_8_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_8_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_8_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_8_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_8_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_8_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_8_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_8_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_8_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_8_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_8_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_8_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_8_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_8_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_9_io_en_r = io_en_a == 7'h9; // @[system.scala 32:27]
  assign rules_9_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_9_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_9_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_9_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_9_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_9_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_9_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_9_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_9_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_9_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_9_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_9_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_9_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_9_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_9_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_9_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_9_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_9_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_10_io_en_r = io_en_a == 7'ha; // @[system.scala 32:27]
  assign rules_10_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_10_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_10_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_10_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_10_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_10_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_10_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_10_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_10_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_10_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_10_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_10_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_10_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_10_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_10_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_10_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_10_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_10_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_11_io_en_r = io_en_a == 7'hb; // @[system.scala 32:27]
  assign rules_11_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_11_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_11_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_11_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_11_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_11_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_11_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_11_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_11_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_11_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_11_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_11_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_11_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_11_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_11_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_11_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_11_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_11_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_12_io_en_r = io_en_a == 7'hc; // @[system.scala 32:27]
  assign rules_12_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_12_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_12_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_12_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_12_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_12_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_12_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_12_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_12_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_12_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_12_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_12_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_12_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_12_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_12_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_12_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_12_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_12_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_13_io_en_r = io_en_a == 7'hd; // @[system.scala 32:27]
  assign rules_13_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_13_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_13_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_13_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_13_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_13_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_13_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_13_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_13_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_13_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_13_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_13_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_13_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_13_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_13_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_13_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_13_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_13_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_14_io_en_r = io_en_a == 7'he; // @[system.scala 32:27]
  assign rules_14_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_14_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_14_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_14_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_14_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_14_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_14_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_14_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_14_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_14_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_14_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_14_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_14_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_14_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_14_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_14_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_14_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_14_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_15_io_en_r = io_en_a == 7'hf; // @[system.scala 32:27]
  assign rules_15_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_15_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_15_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_15_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_15_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_15_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_15_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_15_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_15_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_15_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_15_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_15_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_15_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_15_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_15_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_15_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_15_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_15_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_16_io_en_r = io_en_a == 7'h10; // @[system.scala 32:27]
  assign rules_16_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_16_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_16_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_16_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_16_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_16_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_16_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_16_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_16_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_16_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_16_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_16_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_16_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_16_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_16_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_16_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_16_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_16_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_17_io_en_r = io_en_a == 7'h11; // @[system.scala 32:27]
  assign rules_17_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_17_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_17_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_17_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_17_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_17_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_17_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_17_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_17_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_17_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_17_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_17_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_17_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_17_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_17_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_17_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_17_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_17_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_18_io_en_r = io_en_a == 7'h12; // @[system.scala 32:27]
  assign rules_18_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_18_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_18_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_18_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_18_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_18_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_18_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_18_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_18_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_18_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_18_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_18_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_18_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_18_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_18_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_18_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_18_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_18_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_19_io_en_r = io_en_a == 7'h13; // @[system.scala 32:27]
  assign rules_19_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_19_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_19_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_19_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_19_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_19_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_19_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_19_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_19_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_19_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_19_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_19_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_19_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_19_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_19_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_19_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_19_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_19_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_20_io_en_r = io_en_a == 7'h14; // @[system.scala 32:27]
  assign rules_20_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_20_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_20_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_20_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_20_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_20_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_20_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_20_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_20_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_20_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_20_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_20_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_20_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_20_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_20_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_20_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_20_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_20_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_21_io_en_r = io_en_a == 7'h15; // @[system.scala 32:27]
  assign rules_21_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_21_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_21_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_21_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_21_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_21_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_21_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_21_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_21_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_21_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_21_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_21_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_21_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_21_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_21_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_21_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_21_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_21_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_22_io_en_r = io_en_a == 7'h16; // @[system.scala 32:27]
  assign rules_22_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_22_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_22_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_22_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_22_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_22_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_22_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_22_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_22_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_22_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_22_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_22_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_22_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_22_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_22_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_22_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_22_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_22_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_23_io_en_r = io_en_a == 7'h17; // @[system.scala 32:27]
  assign rules_23_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_23_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_23_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_23_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_23_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_23_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_23_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_23_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_23_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_23_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_23_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_23_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_23_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_23_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_23_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_23_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_23_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_23_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_24_io_en_r = io_en_a == 7'h18; // @[system.scala 32:27]
  assign rules_24_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_24_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_24_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_24_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_24_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_24_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_24_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_24_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_24_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_24_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_24_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_24_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_24_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_24_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_24_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_24_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_24_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_24_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_25_io_en_r = io_en_a == 7'h19; // @[system.scala 32:27]
  assign rules_25_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_25_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_25_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_25_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_25_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_25_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_25_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_25_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_25_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_25_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_25_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_25_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_25_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_25_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_25_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_25_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_25_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_25_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_26_io_en_r = io_en_a == 7'h1a; // @[system.scala 32:27]
  assign rules_26_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_26_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_26_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_26_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_26_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_26_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_26_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_26_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_26_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_26_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_26_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_26_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_26_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_26_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_26_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_26_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_26_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_26_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_27_io_en_r = io_en_a == 7'h1b; // @[system.scala 32:27]
  assign rules_27_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_27_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_27_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_27_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_27_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_27_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_27_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_27_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_27_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_27_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_27_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_27_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_27_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_27_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_27_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_27_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_27_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_27_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_28_io_en_r = io_en_a == 7'h1c; // @[system.scala 32:27]
  assign rules_28_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_28_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_28_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_28_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_28_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_28_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_28_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_28_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_28_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_28_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_28_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_28_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_28_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_28_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_28_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_28_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_28_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_28_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_29_io_en_r = io_en_a == 7'h1d; // @[system.scala 32:27]
  assign rules_29_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_29_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_29_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_29_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_29_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_29_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_29_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_29_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_29_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_29_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_29_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_29_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_29_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_29_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_29_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_29_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_29_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_29_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_30_io_en_r = io_en_a == 7'h1e; // @[system.scala 32:27]
  assign rules_30_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_30_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_30_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_30_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_30_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_30_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_30_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_30_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_30_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_30_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_30_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_30_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_30_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_30_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_30_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_30_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_30_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_30_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_31_io_en_r = io_en_a == 7'h1f; // @[system.scala 32:27]
  assign rules_31_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_31_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_31_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_31_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_31_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_31_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_31_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_31_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_31_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_31_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_31_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_31_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_31_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_31_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_31_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_31_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_31_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_31_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_32_io_en_r = io_en_a == 7'h20; // @[system.scala 32:27]
  assign rules_32_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_32_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_32_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_32_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_32_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_32_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_32_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_32_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_32_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_32_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_32_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_32_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_32_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_32_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_32_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_32_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_32_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_32_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_33_io_en_r = io_en_a == 7'h21; // @[system.scala 32:27]
  assign rules_33_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_33_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_33_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_33_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_33_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_33_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_33_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_33_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_33_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_33_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_33_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_33_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_33_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_33_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_33_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_33_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_33_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_33_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_34_io_en_r = io_en_a == 7'h22; // @[system.scala 32:27]
  assign rules_34_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_34_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_34_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_34_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_34_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_34_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_34_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_34_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_34_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_34_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_34_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_34_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_34_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_34_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_34_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_34_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_34_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_34_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_35_io_en_r = io_en_a == 7'h23; // @[system.scala 32:27]
  assign rules_35_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_35_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_35_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_35_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_35_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_35_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_35_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_35_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_35_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_35_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_35_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_35_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_35_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_35_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_35_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_35_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_35_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_35_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_36_io_en_r = io_en_a == 7'h24; // @[system.scala 32:27]
  assign rules_36_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_36_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_36_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_36_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_36_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_36_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_36_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_36_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_36_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_36_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_36_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_36_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_36_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_36_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_36_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_36_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_36_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_36_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_37_io_en_r = io_en_a == 7'h25; // @[system.scala 32:27]
  assign rules_37_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_37_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_37_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_37_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_37_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_37_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_37_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_37_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_37_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_37_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_37_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_37_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_37_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_37_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_37_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_37_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_37_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_37_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_38_io_en_r = io_en_a == 7'h26; // @[system.scala 32:27]
  assign rules_38_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_38_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_38_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_38_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_38_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_38_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_38_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_38_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_38_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_38_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_38_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_38_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_38_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_38_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_38_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_38_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_38_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_38_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_39_io_en_r = io_en_a == 7'h27; // @[system.scala 32:27]
  assign rules_39_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_39_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_39_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_39_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_39_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_39_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_39_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_39_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_39_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_39_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_39_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_39_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_39_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_39_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_39_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_39_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_39_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_39_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_40_io_en_r = io_en_a == 7'h28; // @[system.scala 32:27]
  assign rules_40_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_40_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_40_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_40_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_40_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_40_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_40_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_40_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_40_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_40_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_40_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_40_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_40_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_40_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_40_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_40_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_40_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_40_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_41_io_en_r = io_en_a == 7'h29; // @[system.scala 32:27]
  assign rules_41_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_41_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_41_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_41_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_41_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_41_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_41_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_41_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_41_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_41_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_41_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_41_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_41_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_41_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_41_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_41_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_41_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_41_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_42_io_en_r = io_en_a == 7'h2a; // @[system.scala 32:27]
  assign rules_42_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_42_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_42_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_42_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_42_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_42_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_42_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_42_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_42_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_42_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_42_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_42_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_42_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_42_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_42_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_42_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_42_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_42_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_43_io_en_r = io_en_a == 7'h2b; // @[system.scala 32:27]
  assign rules_43_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_43_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_43_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_43_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_43_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_43_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_43_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_43_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_43_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_43_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_43_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_43_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_43_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_43_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_43_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_43_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_43_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_43_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_44_io_en_r = io_en_a == 7'h2c; // @[system.scala 32:27]
  assign rules_44_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_44_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_44_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_44_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_44_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_44_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_44_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_44_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_44_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_44_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_44_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_44_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_44_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_44_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_44_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_44_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_44_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_44_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_45_io_en_r = io_en_a == 7'h2d; // @[system.scala 32:27]
  assign rules_45_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_45_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_45_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_45_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_45_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_45_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_45_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_45_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_45_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_45_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_45_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_45_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_45_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_45_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_45_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_45_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_45_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_45_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_46_io_en_r = io_en_a == 7'h2e; // @[system.scala 32:27]
  assign rules_46_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_46_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_46_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_46_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_46_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_46_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_46_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_46_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_46_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_46_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_46_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_46_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_46_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_46_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_46_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_46_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_46_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_46_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_47_io_en_r = io_en_a == 7'h2f; // @[system.scala 32:27]
  assign rules_47_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_47_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_47_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_47_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_47_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_47_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_47_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_47_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_47_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_47_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_47_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_47_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_47_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_47_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_47_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_47_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_47_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_47_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_48_io_en_r = io_en_a == 7'h30; // @[system.scala 32:27]
  assign rules_48_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_48_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_48_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_48_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_48_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_48_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_48_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_48_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_48_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_48_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_48_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_48_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_48_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_48_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_48_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_48_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_48_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_48_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_49_io_en_r = io_en_a == 7'h31; // @[system.scala 32:27]
  assign rules_49_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_49_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_49_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_49_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_49_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_49_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_49_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_49_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_49_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_49_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_49_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_49_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_49_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_49_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_49_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_49_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_49_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_49_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_50_io_en_r = io_en_a == 7'h32; // @[system.scala 32:27]
  assign rules_50_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_50_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_50_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_50_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_50_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_50_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_50_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_50_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_50_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_50_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_50_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_50_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_50_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_50_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_50_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_50_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_50_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_50_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_51_io_en_r = io_en_a == 7'h33; // @[system.scala 32:27]
  assign rules_51_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_51_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_51_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_51_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_51_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_51_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_51_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_51_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_51_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_51_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_51_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_51_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_51_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_51_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_51_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_51_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_51_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_51_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_52_io_en_r = io_en_a == 7'h34; // @[system.scala 32:27]
  assign rules_52_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_52_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_52_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_52_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_52_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_52_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_52_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_52_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_52_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_52_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_52_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_52_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_52_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_52_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_52_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_52_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_52_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_52_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_53_io_en_r = io_en_a == 7'h35; // @[system.scala 32:27]
  assign rules_53_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_53_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_53_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_53_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_53_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_53_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_53_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_53_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_53_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_53_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_53_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_53_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_53_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_53_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_53_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_53_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_53_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_53_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_54_io_en_r = io_en_a == 7'h36; // @[system.scala 32:27]
  assign rules_54_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_54_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_54_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_54_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_54_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_54_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_54_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_54_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_54_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_54_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_54_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_54_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_54_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_54_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_54_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_54_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_54_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_54_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_55_io_en_r = io_en_a == 7'h37; // @[system.scala 32:27]
  assign rules_55_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_55_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_55_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_55_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_55_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_55_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_55_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_55_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_55_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_55_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_55_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_55_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_55_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_55_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_55_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_55_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_55_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_55_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_56_io_en_r = io_en_a == 7'h38; // @[system.scala 32:27]
  assign rules_56_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_56_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_56_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_56_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_56_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_56_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_56_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_56_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_56_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_56_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_56_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_56_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_56_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_56_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_56_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_56_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_56_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_56_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_57_io_en_r = io_en_a == 7'h39; // @[system.scala 32:27]
  assign rules_57_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_57_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_57_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_57_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_57_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_57_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_57_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_57_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_57_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_57_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_57_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_57_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_57_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_57_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_57_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_57_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_57_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_57_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_58_io_en_r = io_en_a == 7'h3a; // @[system.scala 32:27]
  assign rules_58_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_58_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_58_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_58_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_58_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_58_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_58_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_58_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_58_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_58_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_58_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_58_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_58_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_58_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_58_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_58_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_58_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_58_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_59_io_en_r = io_en_a == 7'h3b; // @[system.scala 32:27]
  assign rules_59_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_59_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_59_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_59_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_59_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_59_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_59_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_59_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_59_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_59_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_59_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_59_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_59_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_59_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_59_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_59_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_59_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_59_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_60_io_en_r = io_en_a == 7'h3c; // @[system.scala 32:27]
  assign rules_60_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_60_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_60_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_60_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_60_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_60_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_60_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_60_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_60_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_60_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_60_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_60_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_60_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_60_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_60_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_60_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_60_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_60_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_61_io_en_r = io_en_a == 7'h3d; // @[system.scala 32:27]
  assign rules_61_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_61_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_61_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_61_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_61_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_61_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_61_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_61_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_61_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_61_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_61_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_61_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_61_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_61_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_61_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_61_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_61_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_61_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_62_io_en_r = io_en_a == 7'h3e; // @[system.scala 32:27]
  assign rules_62_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_62_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_62_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_62_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_62_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_62_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_62_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_62_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_62_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_62_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_62_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_62_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_62_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_62_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_62_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_62_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_62_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_62_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_63_io_en_r = io_en_a == 7'h3f; // @[system.scala 32:27]
  assign rules_63_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_63_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_63_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_63_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_63_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_63_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_63_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_63_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_63_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_63_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_63_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_63_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_63_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_63_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_63_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_63_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_63_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_63_io_x_in = x_reg; // @[system.scala 31:18]
  assign rules_64_io_en_r = io_en_a == 7'h40; // @[system.scala 32:27]
  assign rules_64_io_n_in_0 = n_reg_0; // @[system.scala 30:18]
  assign rules_64_io_n_in_1 = n_reg_1; // @[system.scala 30:18]
  assign rules_64_io_n_in_2 = n_reg_2; // @[system.scala 30:18]
  assign rules_64_io_n_in_3 = n_reg_3; // @[system.scala 30:18]
  assign rules_64_io_n_in_4 = n_reg_4; // @[system.scala 30:18]
  assign rules_64_io_n_in_5 = n_reg_5; // @[system.scala 30:18]
  assign rules_64_io_n_in_6 = n_reg_6; // @[system.scala 30:18]
  assign rules_64_io_n_in_7 = n_reg_7; // @[system.scala 30:18]
  assign rules_64_io_n_in_8 = n_reg_8; // @[system.scala 30:18]
  assign rules_64_io_n_in_9 = n_reg_9; // @[system.scala 30:18]
  assign rules_64_io_n_in_10 = n_reg_10; // @[system.scala 30:18]
  assign rules_64_io_n_in_11 = n_reg_11; // @[system.scala 30:18]
  assign rules_64_io_n_in_12 = n_reg_12; // @[system.scala 30:18]
  assign rules_64_io_n_in_13 = n_reg_13; // @[system.scala 30:18]
  assign rules_64_io_n_in_14 = n_reg_14; // @[system.scala 30:18]
  assign rules_64_io_n_in_15 = n_reg_15; // @[system.scala 30:18]
  assign rules_64_io_n_in_16 = n_reg_16; // @[system.scala 30:18]
  assign rules_64_io_x_in = x_reg; // @[system.scala 31:18]
  always @(posedge clock) begin
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_0 <= rules_64_io_n_out_0; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_0 <= rules_63_io_n_out_0; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_0 <= rules_62_io_n_out_0; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_0 <= rules_61_io_n_out_0; // @[system.scala 34:7]
    end else begin
      n_reg_0 <= _GEN_1080;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_1 <= rules_64_io_n_out_1; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_1 <= rules_63_io_n_out_1; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_1 <= rules_62_io_n_out_1; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_1 <= rules_61_io_n_out_1; // @[system.scala 34:7]
    end else begin
      n_reg_1 <= _GEN_1081;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_2 <= rules_64_io_n_out_2; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_2 <= rules_63_io_n_out_2; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_2 <= rules_62_io_n_out_2; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_2 <= rules_61_io_n_out_2; // @[system.scala 34:7]
    end else begin
      n_reg_2 <= _GEN_1082;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_3 <= rules_64_io_n_out_3; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_3 <= rules_63_io_n_out_3; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_3 <= rules_62_io_n_out_3; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_3 <= rules_61_io_n_out_3; // @[system.scala 34:7]
    end else begin
      n_reg_3 <= _GEN_1083;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_4 <= rules_64_io_n_out_4; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_4 <= rules_63_io_n_out_4; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_4 <= rules_62_io_n_out_4; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_4 <= rules_61_io_n_out_4; // @[system.scala 34:7]
    end else begin
      n_reg_4 <= _GEN_1084;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_5 <= rules_64_io_n_out_5; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_5 <= rules_63_io_n_out_5; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_5 <= rules_62_io_n_out_5; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_5 <= rules_61_io_n_out_5; // @[system.scala 34:7]
    end else begin
      n_reg_5 <= _GEN_1085;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_6 <= rules_64_io_n_out_6; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_6 <= rules_63_io_n_out_6; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_6 <= rules_62_io_n_out_6; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_6 <= rules_61_io_n_out_6; // @[system.scala 34:7]
    end else begin
      n_reg_6 <= _GEN_1086;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_7 <= rules_64_io_n_out_7; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_7 <= rules_63_io_n_out_7; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_7 <= rules_62_io_n_out_7; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_7 <= rules_61_io_n_out_7; // @[system.scala 34:7]
    end else begin
      n_reg_7 <= _GEN_1087;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_8 <= rules_64_io_n_out_8; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_8 <= rules_63_io_n_out_8; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_8 <= rules_62_io_n_out_8; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_8 <= rules_61_io_n_out_8; // @[system.scala 34:7]
    end else begin
      n_reg_8 <= _GEN_1088;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_9 <= rules_64_io_n_out_9; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_9 <= rules_63_io_n_out_9; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_9 <= rules_62_io_n_out_9; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_9 <= rules_61_io_n_out_9; // @[system.scala 34:7]
    end else begin
      n_reg_9 <= _GEN_1089;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_10 <= rules_64_io_n_out_10; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_10 <= rules_63_io_n_out_10; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_10 <= rules_62_io_n_out_10; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_10 <= rules_61_io_n_out_10; // @[system.scala 34:7]
    end else begin
      n_reg_10 <= _GEN_1090;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_11 <= rules_64_io_n_out_11; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_11 <= rules_63_io_n_out_11; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_11 <= rules_62_io_n_out_11; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_11 <= rules_61_io_n_out_11; // @[system.scala 34:7]
    end else begin
      n_reg_11 <= _GEN_1091;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_12 <= rules_64_io_n_out_12; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_12 <= rules_63_io_n_out_12; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_12 <= rules_62_io_n_out_12; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_12 <= rules_61_io_n_out_12; // @[system.scala 34:7]
    end else begin
      n_reg_12 <= _GEN_1092;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_13 <= rules_64_io_n_out_13; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_13 <= rules_63_io_n_out_13; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_13 <= rules_62_io_n_out_13; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_13 <= rules_61_io_n_out_13; // @[system.scala 34:7]
    end else begin
      n_reg_13 <= _GEN_1093;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_14 <= rules_64_io_n_out_14; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_14 <= rules_63_io_n_out_14; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_14 <= rules_62_io_n_out_14; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_14 <= rules_61_io_n_out_14; // @[system.scala 34:7]
    end else begin
      n_reg_14 <= _GEN_1094;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_15 <= rules_64_io_n_out_15; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_15 <= rules_63_io_n_out_15; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_15 <= rules_62_io_n_out_15; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_15 <= rules_61_io_n_out_15; // @[system.scala 34:7]
    end else begin
      n_reg_15 <= _GEN_1095;
    end
    if (_T_128) begin // @[system.scala 33:21]
      n_reg_16 <= rules_64_io_n_out_16; // @[system.scala 34:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      n_reg_16 <= rules_63_io_n_out_16; // @[system.scala 34:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      n_reg_16 <= rules_62_io_n_out_16; // @[system.scala 34:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      n_reg_16 <= rules_61_io_n_out_16; // @[system.scala 34:7]
    end else begin
      n_reg_16 <= _GEN_1096;
    end
    if (_T_128) begin // @[system.scala 33:21]
      x_reg <= rules_64_io_x_out; // @[system.scala 35:7]
    end else if (_T_126) begin // @[system.scala 33:21]
      x_reg <= rules_63_io_x_out; // @[system.scala 35:7]
    end else if (_T_124) begin // @[system.scala 33:21]
      x_reg <= rules_62_io_x_out; // @[system.scala 35:7]
    end else if (_T_122) begin // @[system.scala 33:21]
      x_reg <= rules_61_io_x_out; // @[system.scala 35:7]
    end else begin
      x_reg <= _GEN_1097;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif

                initial begin
                    assume(reset==1 && io_en_a==0);
                end

                  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_1 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_2 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_3 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_4 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_5 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_6 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_7 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_8 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_9 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_10 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_11 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_12 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_13 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_14 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_15 == 2'h2) | n_reg_16 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_1 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_2 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_3 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_4 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_5 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_6 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_7 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_8 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_9 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_10 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_11 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_12 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_13 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_14 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(~(n_reg_16 == 2'h2) | n_reg_15 != 2'h2); // @[system.scala 57:7]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[system.scala 57:7]
    end
  end
endmodule
